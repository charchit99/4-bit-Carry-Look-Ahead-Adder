magic
tech scmos
timestamp 1618889747
<< nwell >>
rect -19 -3 5 17
<< ntransistor >>
rect -8 -13 -6 -9
<< ptransistor >>
rect -8 3 -6 11
<< ndiffusion >>
rect -9 -13 -8 -9
rect -6 -13 -5 -9
<< pdiffusion >>
rect -9 3 -8 11
rect -6 3 -5 11
<< ndcontact >>
rect -13 -13 -9 -9
rect -5 -13 -1 -9
<< pdcontact >>
rect -13 3 -9 11
rect -5 3 -1 11
<< polysilicon >>
rect -8 11 -6 14
rect -8 -9 -6 3
rect -8 -16 -6 -13
<< polycontact >>
rect -12 -6 -8 -2
<< metal1 >>
rect -19 15 5 18
rect -13 11 -9 15
rect -5 -2 -1 3
rect -19 -6 -12 -2
rect -5 -6 5 -2
rect -5 -9 -1 -6
rect -13 -17 -9 -13
rect -19 -20 5 -17
<< labels >>
rlabel metal1 -13 17 -2 18 5 vdd
rlabel metal1 -19 -4 -15 -3 3 input
rlabel metal1 1 -4 5 -3 7 output
rlabel metal1 -9 -20 -5 -19 1 gnd
<< end >>

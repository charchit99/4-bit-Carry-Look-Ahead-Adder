* SPICE3 file created from sum.ext - technology: scmos

.option scale=0.09u

M1000 xs10 c1_bar vdd w_12_n49# pfet w=8 l=2
+  ad=48 pd=28 as=640 ps=416
M1001 s1 p1 xs10 w_12_n49# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1002 xs30 c3_bar vdd w_170_n49# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 s3 p3 xs30 w_170_n49# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1004 xs11 c1 vdd w_12_n49# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1005 s1 p1_bar xs11 w_12_n49# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 xs31 c3 vdd w_170_n49# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1007 s3 p3_bar xs31 w_170_n49# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 c1_bar c1 vdd w_n58_n60# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1009 p1_bar p1 vdd w_n58_n60# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1010 c3_bar c3 vdd w_100_n60# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1011 p3_bar p3 vdd w_100_n60# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1012 c1_bar c1 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=320 ps=288
M1013 p1_bar p1 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1014 xs12 c1 gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1015 s1 p1 xs12 Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1016 c3_bar c3 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 p3_bar p3 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 xs32 c3 gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1019 s3 p3 xs32 Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1020 xs13 c1_bar gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1021 s1 p1_bar xs13 Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 xs33 c3_bar gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1023 s3 p3_bar xs33 Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 xs00 c0_bar vdd w_12_n147# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1025 s0 p0 xs00 w_12_n147# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1026 xs20 c2_bar vdd w_170_n147# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1027 s2 p2 xs20 w_170_n147# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1028 xs01 c0 vdd w_12_n147# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1029 s0 p0_bar xs01 w_12_n147# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 xs21 c2 vdd w_170_n147# pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1031 s2 p2_bar xs21 w_170_n147# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 c0_bar c0 vdd w_n58_n158# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1033 p0_bar p0 vdd w_n58_n158# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1034 c2_bar c2 vdd w_100_n158# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1035 p2_bar p2 vdd w_100_n158# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1036 c0_bar c0 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1037 p0_bar p0 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1038 xs02 c0 gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1039 s0 p0 xs02 Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1040 c2_bar c2 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1041 p2_bar p2 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1042 xs22 c2 gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1043 s2 p2 xs22 Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1044 xs03 c0_bar gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1045 s0 p0_bar xs03 Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 xs23 c2_bar gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1047 s2 p2_bar xs23 Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 c0 gnd 0.86fF
C1 vdd c0_bar 0.48fF
C2 p1 p2 0.34fF
C3 c1 gnd 0.77fF
C4 s1 xs13 0.04fF
C5 p0_bar vdd 0.17fF
C6 s2 s1 0.25fF
C7 w_n58_n158# c0_bar 0.08fF
C8 p3 c3 0.23fF
C9 vdd p1_bar 0.25fF
C10 s1 s3 0.09fF
C11 c3_bar p3_bar 0.12fF
C12 w_n58_n158# p0_bar 0.16fF
C13 w_12_n147# c0 0.06fF
C14 w_170_n49# c3 0.06fF
C15 w_12_n49# xs11 0.01fF
C16 w_100_n60# p3_bar 0.16fF
C17 c1_bar vdd 0.44fF
C18 s2 xs20 0.08fF
C19 w_100_n60# c3_bar 0.08fF
C20 w_n58_n60# vdd 0.11fF
C21 vdd s0 1.32fF
C22 w_12_n147# xs00 0.01fF
C23 c2_bar p2 0.04fF
C24 p2_bar p2 0.37fF
C25 gnd c0_bar 0.18fF
C26 p0_bar gnd 0.04fF
C27 s3 xs32 0.04fF
C28 vdd p0 0.34fF
C29 p1_bar gnd 0.04fF
C30 c2 vdd 0.04fF
C31 w_12_n147# c0_bar 0.19fF
C32 w_n58_n158# p0 0.14fF
C33 p3 p3_bar 0.37fF
C34 vdd c3 0.17fF
C35 xs30 s3 0.08fF
C36 c1_bar gnd 0.18fF
C37 w_12_n147# p0_bar 0.29fF
C38 xs02 s0 0.04fF
C39 w_170_n49# p3_bar 0.27fF
C40 c3_bar p3 0.04fF
C41 p1 vdd 0.16fF
C42 w_12_n49# vdd 0.06fF
C43 w_170_n49# c3_bar 0.19fF
C44 w_100_n60# p3 0.14fF
C45 w_12_n147# s0 0.06fF
C46 w_170_n147# xs20 0.01fF
C47 s2 xs23 0.04fF
C48 gnd p0 0.33fF
C49 c2 gnd 1.83fF
C50 p3 p2 1.58fF
C51 vdd c2_bar 0.48fF
C52 c3 gnd 0.68fF
C53 p2_bar vdd 0.17fF
C54 s2 s3 0.59fF
C55 w_12_n147# p0 0.19fF
C56 s1 p1_bar 0.46fF
C57 p1 gnd 0.14fF
C58 vdd p3_bar 0.25fF
C59 c3_bar vdd 0.44fF
C60 w_12_n49# xs10 0.01fF
C61 w_100_n60# vdd 0.11fF
C62 w_170_n49# p3 0.19fF
C63 s1 s0 1.25fF
C64 gnd c2_bar 0.18fF
C65 p2_bar gnd 0.04fF
C66 p3_bar gnd 0.04fF
C67 vdd p2 1.35fF
C68 s3 xs33 0.04fF
C69 xs01 vdd 0.08fF
C70 vdd xs11 0.08fF
C71 c3_bar gnd 0.18fF
C72 xs03 s0 0.04fF
C73 s2 w_170_n147# 0.06fF
C74 w_170_n49# xs31 0.01fF
C75 p3 vdd 0.16fF
C76 p1 s1 0.45fF
C77 w_170_n49# vdd 0.06fF
C78 w_12_n49# s1 0.06fF
C79 gnd p2 0.33fF
C80 xs21 vdd 0.08fF
C81 c0 c1 0.19fF
C82 p3 gnd 0.14fF
C83 vdd xs31 0.08fF
C84 w_12_n147# xs01 0.01fF
C85 s2 s0 0.09fF
C86 w_n58_n158# vdd 0.11fF
C87 s3 s0 0.09fF
C88 c0 c0_bar 0.16fF
C89 s1 p2 0.07fF
C90 c0 p0_bar 0.04fF
C91 c1 p1_bar 0.04fF
C92 vdd gnd 0.39fF
C93 s1 xs11 0.08fF
C94 c2 w_100_n158# 0.11fF
C95 c1_bar c1 0.16fF
C96 p3 s1 0.07fF
C97 vdd xs10 0.08fF
C98 w_n58_n60# c1 0.11fF
C99 w_12_n147# vdd 0.06fF
C100 xs00 s0 0.08fF
C101 xs02 gnd 0.04fF
C102 c0 p0 0.24fF
C103 p0_bar c0_bar 0.12fF
C104 c0 c2 0.05fF
C105 s2 p2_bar 0.45fF
C106 c1 p0 0.07fF
C107 c2 c1 0.09fF
C108 s3 p3_bar 0.45fF
C109 w_100_n158# c2_bar 0.08fF
C110 p2_bar w_100_n158# 0.16fF
C111 c2 w_170_n147# 0.06fF
C112 c1_bar p1_bar 0.12fF
C113 p1 c1 0.23fF
C114 vdd s1 0.35fF
C115 p0_bar s0 0.53fF
C116 w_n58_n60# p1_bar 0.16fF
C117 w_170_n49# xs30 0.01fF
C118 w_12_n49# c1 0.06fF
C119 p1_bar s0 0.10fF
C120 w_n58_n60# c1_bar 0.08fF
C121 vdd xs20 0.08fF
C122 c0_bar p0 0.04fF
C123 xs22 gnd 0.04fF
C124 s2 p2 0.45fF
C125 p0_bar p0 0.37fF
C126 gnd xs12 0.04fF
C127 w_100_n158# p2 0.14fF
C128 w_170_n147# c2_bar 0.19fF
C129 p2_bar w_170_n147# 0.29fF
C130 p0 s0 0.45fF
C131 p1 p1_bar 0.37fF
C132 p3 s3 0.45fF
C133 xs10 s1 0.08fF
C134 vdd xs30 0.08fF
C135 w_170_n49# s3 0.06fF
C136 w_12_n49# p1_bar 0.27fF
C137 c3 s0 0.19fF
C138 c1_bar p1 0.04fF
C139 w_n58_n60# p1 0.14fF
C140 w_12_n49# c1_bar 0.19fF
C141 xs03 gnd 0.04fF
C142 gnd xs32 0.04fF
C143 s2 xs21 0.08fF
C144 c2 c3 1.57fF
C145 s1 xs12 0.04fF
C146 s3 xs31 0.08fF
C147 w_170_n147# p2 0.19fF
C148 p1 p0 0.13fF
C149 s2 vdd 0.11fF
C150 vdd s3 0.11fF
C151 w_100_n158# vdd 0.11fF
C152 w_12_n49# p1 0.19fF
C153 c2 c2_bar 0.16fF
C154 xs23 gnd 0.04fF
C155 c2 p2_bar 0.04fF
C156 gnd xs13 0.04fF
C157 c3 p3_bar 0.04fF
C158 c0 vdd 0.04fF
C159 xs21 w_170_n147# 0.01fF
C160 p2 s0 0.07fF
C161 vdd c1 0.17fF
C162 c3_bar c3 0.16fF
C163 w_n58_n158# c0 0.11fF
C164 xs01 s0 0.08fF
C165 w_100_n60# c3 0.11fF
C166 w_170_n147# vdd 0.06fF
C167 vdd xs00 0.08fF
C168 p3 s0 0.07fF
C169 c2 p2 0.24fF
C170 p2_bar c2_bar 0.12fF
C171 gnd xs33 0.04fF
C172 c3 p2 0.07fF
C173 s2 xs22 0.04fF
C174 xs23 Gnd 0.01fF
C175 xs03 Gnd 0.01fF
C176 xs22 Gnd 0.01fF
C177 xs02 Gnd 0.01fF
C178 xs21 Gnd 0.00fF
C179 xs01 Gnd 0.00fF
C180 p2_bar Gnd 0.02fF
C181 c2 Gnd 2.56fF
C182 p0_bar Gnd 0.02fF
C183 c0 Gnd 1.98fF
C184 s2 Gnd 1.41fF
C185 xs20 Gnd 0.00fF
C186 s0 Gnd 3.27fF
C187 xs00 Gnd 0.00fF
C188 p2 Gnd 1.59fF
C189 c2_bar Gnd 0.42fF
C190 p0 Gnd 1.02fF
C191 c0_bar Gnd 0.02fF
C192 xs33 Gnd 0.01fF
C193 xs13 Gnd 0.01fF
C194 xs32 Gnd 0.01fF
C195 xs12 Gnd 0.01fF
C196 gnd Gnd 1.16fF
C197 xs31 Gnd 0.00fF
C198 xs11 Gnd 0.00fF
C199 p3_bar Gnd 0.21fF
C200 c3 Gnd 3.80fF
C201 p1_bar Gnd 2.16fF
C202 c1 Gnd 3.26fF
C203 s3 Gnd 1.17fF
C204 xs30 Gnd 0.00fF
C205 s1 Gnd 1.75fF
C206 xs10 Gnd 0.00fF
C207 vdd Gnd 3.49fF
C208 p3 Gnd 0.23fF
C209 c3_bar Gnd 0.42fF
C210 p1 Gnd 1.01fF
C211 c1_bar Gnd 0.42fF
C212 w_170_n147# Gnd 1.35fF
C213 w_100_n158# Gnd 1.08fF
C214 w_12_n147# Gnd 1.35fF
C215 w_n58_n158# Gnd 1.08fF
C216 w_170_n49# Gnd 0.13fF
C217 w_100_n60# Gnd 1.08fF
C218 w_12_n49# Gnd 1.35fF
C219 w_n58_n60# Gnd 1.08fF

magic
tech scmos
timestamp 1619396629
<< nwell >>
rect -49 23 39 43
rect 106 23 172 43
rect 225 23 271 43
rect 326 25 352 45
rect -39 -14 29 6
rect 116 -14 172 6
rect 235 -7 282 13
rect 326 -1 362 19
rect 362 -50 388 -30
rect 281 -74 308 -54
rect 41 -116 68 -96
rect 176 -98 203 -78
<< ntransistor >>
rect 338 -35 340 -31
rect 348 -35 350 -31
rect 247 -58 249 -54
rect 257 -58 259 -54
rect 267 -58 269 -54
rect 338 -58 340 -54
rect 374 -60 376 -56
rect 128 -82 130 -78
rect 138 -82 140 -78
rect 148 -82 150 -78
rect 158 -82 160 -78
rect 247 -85 249 -81
rect 267 -85 269 -81
rect 293 -85 295 -81
rect -27 -100 -25 -96
rect -17 -100 -15 -96
rect -7 -100 -5 -96
rect 3 -100 5 -96
rect 13 -100 15 -96
rect 128 -109 130 -105
rect 148 -109 150 -105
rect 168 -109 170 -105
rect 188 -109 190 -105
rect -27 -127 -25 -123
rect -7 -127 -5 -123
rect 13 -127 15 -123
rect 33 -127 35 -123
rect 53 -127 55 -123
<< ptransistor >>
rect -37 29 -35 37
rect -17 29 -15 37
rect 3 29 5 37
rect 23 29 25 37
rect 118 29 120 37
rect 138 29 140 37
rect 158 29 160 37
rect 237 29 239 37
rect 257 29 259 37
rect 338 31 340 39
rect -27 -8 -25 0
rect -17 -8 -15 0
rect -7 -8 -5 0
rect 3 -8 5 0
rect 13 -8 15 0
rect 128 -8 130 0
rect 138 -8 140 0
rect 148 -8 150 0
rect 158 -8 160 0
rect 247 -1 249 7
rect 257 -1 259 7
rect 267 -1 269 7
rect 338 5 340 13
rect 348 5 350 13
rect 374 -44 376 -36
rect 293 -68 295 -60
rect 188 -92 190 -84
rect 53 -110 55 -102
<< ndiffusion >>
rect 336 -35 338 -31
rect 340 -35 342 -31
rect 346 -35 348 -31
rect 350 -35 352 -31
rect 245 -58 247 -54
rect 249 -58 251 -54
rect 255 -58 257 -54
rect 259 -58 261 -54
rect 265 -58 267 -54
rect 269 -58 271 -54
rect 336 -58 338 -54
rect 340 -58 342 -54
rect 372 -60 374 -56
rect 376 -60 378 -56
rect 126 -82 128 -78
rect 130 -82 132 -78
rect 136 -82 138 -78
rect 140 -82 142 -78
rect 146 -82 148 -78
rect 150 -82 152 -78
rect 156 -82 158 -78
rect 160 -82 162 -78
rect 245 -85 247 -81
rect 249 -85 251 -81
rect 265 -85 267 -81
rect 269 -85 271 -81
rect 291 -85 293 -81
rect 295 -85 297 -81
rect -29 -100 -27 -96
rect -25 -100 -23 -96
rect -19 -100 -17 -96
rect -15 -100 -13 -96
rect -9 -100 -7 -96
rect -5 -100 -3 -96
rect 1 -100 3 -96
rect 5 -100 7 -96
rect 11 -100 13 -96
rect 15 -100 17 -96
rect 126 -109 128 -105
rect 130 -109 132 -105
rect 146 -109 148 -105
rect 150 -109 152 -105
rect 166 -109 168 -105
rect 170 -109 172 -105
rect 186 -109 188 -105
rect 190 -109 192 -105
rect -29 -127 -27 -123
rect -25 -127 -23 -123
rect -9 -127 -7 -123
rect -5 -127 -3 -123
rect 11 -127 13 -123
rect 15 -127 17 -123
rect 31 -127 33 -123
rect 35 -127 37 -123
rect 51 -127 53 -123
rect 55 -127 57 -123
<< pdiffusion >>
rect -39 29 -37 37
rect -35 29 -33 37
rect -19 29 -17 37
rect -15 29 -13 37
rect 1 29 3 37
rect 5 29 7 37
rect 21 29 23 37
rect 25 29 27 37
rect 116 29 118 37
rect 120 29 122 37
rect 136 29 138 37
rect 140 29 142 37
rect 156 29 158 37
rect 160 29 162 37
rect 235 29 237 37
rect 239 29 241 37
rect 255 29 257 37
rect 259 29 261 37
rect 336 31 338 39
rect 340 31 342 39
rect -29 -8 -27 0
rect -25 -8 -23 0
rect -19 -8 -17 0
rect -15 -8 -13 0
rect -9 -8 -7 0
rect -5 -8 -3 0
rect 1 -8 3 0
rect 5 -8 7 0
rect 11 -8 13 0
rect 15 -8 17 0
rect 126 -8 128 0
rect 130 -8 132 0
rect 136 -8 138 0
rect 140 -8 142 0
rect 146 -8 148 0
rect 150 -8 152 0
rect 156 -8 158 0
rect 160 -8 162 0
rect 245 -1 247 7
rect 249 -1 251 7
rect 255 -1 257 7
rect 259 -1 261 7
rect 265 -1 267 7
rect 269 -1 271 7
rect 336 5 338 13
rect 340 5 342 13
rect 346 5 348 13
rect 350 5 352 13
rect 372 -44 374 -36
rect 376 -44 378 -36
rect 291 -68 293 -60
rect 295 -68 297 -60
rect 186 -92 188 -84
rect 190 -92 192 -84
rect 51 -110 53 -102
rect 55 -110 57 -102
<< ndcontact >>
rect 332 -35 336 -31
rect 342 -35 346 -31
rect 352 -35 356 -31
rect 241 -58 245 -54
rect 251 -58 255 -54
rect 261 -58 265 -54
rect 271 -58 275 -54
rect 332 -58 336 -54
rect 342 -58 346 -54
rect 368 -60 372 -56
rect 378 -60 382 -56
rect 122 -82 126 -78
rect 132 -82 136 -78
rect 142 -82 146 -78
rect 152 -82 156 -78
rect 162 -82 166 -78
rect 241 -85 245 -81
rect 251 -85 255 -81
rect 261 -85 265 -81
rect 271 -85 275 -81
rect 287 -85 291 -81
rect 297 -85 301 -81
rect -33 -100 -29 -96
rect -23 -100 -19 -96
rect -13 -100 -9 -96
rect -3 -100 1 -96
rect 7 -100 11 -96
rect 17 -100 21 -96
rect 122 -109 126 -105
rect 132 -109 136 -105
rect 142 -109 146 -105
rect 152 -109 156 -105
rect 162 -109 166 -105
rect 172 -109 176 -105
rect 182 -109 186 -105
rect 192 -109 196 -105
rect -33 -127 -29 -123
rect -23 -127 -19 -123
rect -13 -127 -9 -123
rect -3 -127 1 -123
rect 7 -127 11 -123
rect 17 -127 21 -123
rect 27 -127 31 -123
rect 37 -127 41 -123
rect 47 -127 51 -123
rect 57 -127 61 -123
<< pdcontact >>
rect -43 29 -39 37
rect -33 29 -29 37
rect -23 29 -19 37
rect -13 29 -9 37
rect -3 29 1 37
rect 7 29 11 37
rect 17 29 21 37
rect 27 29 31 37
rect 112 29 116 37
rect 122 29 126 37
rect 132 29 136 37
rect 142 29 146 37
rect 152 29 156 37
rect 162 29 166 37
rect 231 29 235 37
rect 241 29 245 37
rect 251 29 255 37
rect 261 29 265 37
rect 332 31 336 39
rect 342 31 346 39
rect -33 -8 -29 0
rect -23 -8 -19 0
rect -13 -8 -9 0
rect -3 -8 1 0
rect 7 -8 11 0
rect 17 -8 21 0
rect 122 -8 126 0
rect 132 -8 136 0
rect 142 -8 146 0
rect 152 -8 156 0
rect 162 -8 166 0
rect 241 -1 245 7
rect 251 -1 255 7
rect 261 -1 265 7
rect 271 -1 275 7
rect 332 5 336 13
rect 342 5 346 13
rect 352 5 356 13
rect 368 -44 372 -36
rect 378 -44 382 -36
rect 287 -68 291 -60
rect 297 -68 301 -60
rect 182 -92 186 -84
rect 192 -92 196 -84
rect 47 -110 51 -102
rect 57 -110 61 -102
<< polysilicon >>
rect -37 37 -35 71
rect -17 37 -15 62
rect 3 37 5 53
rect 23 37 25 44
rect 118 37 120 62
rect 138 37 140 53
rect 158 37 160 44
rect 237 37 239 53
rect 257 37 259 44
rect 338 39 340 46
rect -37 26 -35 29
rect -17 26 -15 29
rect 3 26 5 29
rect 23 26 25 29
rect 118 26 120 29
rect 138 26 140 29
rect 158 26 160 29
rect 237 26 239 29
rect 257 26 259 29
rect 338 28 340 31
rect 338 13 340 16
rect 348 13 350 16
rect 247 7 249 10
rect 257 7 259 10
rect 267 7 269 10
rect -27 0 -25 3
rect -17 0 -15 3
rect -7 0 -5 3
rect 3 0 5 3
rect 13 0 15 3
rect 128 0 130 3
rect 138 0 140 3
rect 148 0 150 3
rect 158 0 160 3
rect -27 -96 -25 -8
rect -17 -15 -15 -8
rect -7 -24 -5 -8
rect 3 -33 5 -8
rect 13 -42 15 -8
rect -17 -96 -15 -62
rect -7 -96 -5 -71
rect 128 -78 130 -8
rect 138 -15 140 -8
rect 148 -24 150 -8
rect 158 -33 160 -8
rect 138 -78 140 -53
rect 247 -54 249 -1
rect 257 -8 259 -1
rect 267 -17 269 -1
rect 338 -31 340 5
rect 348 -2 350 5
rect 348 -31 350 -24
rect 338 -38 340 -35
rect 348 -38 350 -35
rect 374 -36 376 -33
rect 257 -54 259 -38
rect 267 -54 269 -47
rect 338 -54 340 -51
rect 247 -61 249 -58
rect 257 -61 259 -58
rect 267 -61 269 -58
rect 293 -60 295 -57
rect 374 -56 376 -44
rect 148 -78 150 -62
rect 338 -65 340 -58
rect 374 -63 376 -60
rect 158 -78 160 -71
rect 3 -96 5 -80
rect 247 -81 249 -78
rect 267 -81 269 -78
rect 293 -81 295 -68
rect 128 -85 130 -82
rect 138 -85 140 -82
rect 148 -85 150 -82
rect 158 -85 160 -82
rect 188 -84 190 -81
rect 13 -96 15 -89
rect 247 -92 249 -85
rect -27 -103 -25 -100
rect -17 -103 -15 -100
rect -7 -103 -5 -100
rect 3 -103 5 -100
rect 13 -103 15 -100
rect 53 -102 55 -99
rect 128 -105 130 -102
rect 148 -105 150 -102
rect 168 -105 170 -102
rect 188 -105 190 -92
rect 267 -101 269 -85
rect 293 -88 295 -85
rect -27 -123 -25 -120
rect -7 -123 -5 -120
rect 13 -123 15 -120
rect 33 -123 35 -120
rect 53 -123 55 -110
rect 128 -116 130 -109
rect 148 -125 150 -109
rect -27 -134 -25 -127
rect -7 -143 -5 -127
rect 13 -152 15 -127
rect 33 -161 35 -127
rect 53 -130 55 -127
rect 168 -134 170 -109
rect 188 -112 190 -109
<< polycontact >>
rect -35 67 -31 71
rect -15 58 -11 62
rect 5 49 9 53
rect 25 40 29 44
rect 120 58 124 62
rect 140 49 144 53
rect 160 40 164 44
rect 239 49 243 53
rect 259 40 263 44
rect 340 42 344 46
rect -31 -54 -27 -50
rect -21 -15 -17 -11
rect -11 -24 -7 -20
rect -1 -33 3 -29
rect 9 -42 13 -38
rect 124 -46 128 -42
rect -21 -66 -17 -62
rect -11 -75 -7 -71
rect 134 -15 138 -11
rect 144 -24 148 -20
rect 154 -33 158 -29
rect 243 -30 247 -26
rect 134 -57 138 -53
rect 253 -8 257 -4
rect 263 -17 267 -13
rect 334 -15 338 -11
rect 344 -2 348 2
rect 344 -28 348 -24
rect 253 -42 257 -38
rect 263 -51 267 -47
rect 370 -52 374 -48
rect 144 -66 148 -62
rect 334 -65 338 -61
rect 154 -75 158 -71
rect 289 -76 293 -72
rect -1 -84 3 -80
rect 9 -93 13 -89
rect 243 -92 247 -88
rect 184 -100 188 -96
rect 263 -101 267 -97
rect 49 -118 53 -114
rect 124 -116 128 -112
rect 144 -125 148 -121
rect -31 -134 -27 -130
rect -11 -143 -7 -139
rect 9 -152 13 -148
rect 29 -161 33 -157
rect 164 -134 168 -130
<< metal1 >>
rect -31 67 44 71
rect -11 58 -7 62
rect 9 49 13 53
rect 29 40 32 44
rect -43 25 -39 29
rect -43 0 -39 20
rect -33 10 -29 29
rect -23 25 -19 29
rect -33 6 -19 10
rect -23 0 -19 6
rect -43 -4 -33 0
rect -13 0 -9 29
rect -3 25 1 29
rect 7 17 11 29
rect 17 25 21 29
rect -3 13 11 17
rect -3 0 1 13
rect 27 10 31 29
rect 7 6 31 10
rect 7 0 11 6
rect -73 -19 -17 -15
rect -73 -129 -69 -19
rect -65 -28 -7 -24
rect -65 -138 -61 -28
rect -57 -37 3 -33
rect -57 -147 -53 -37
rect -49 -46 13 -42
rect -49 -157 -45 -46
rect 17 -49 21 -8
rect -35 -54 -31 -50
rect 40 -57 44 67
rect 124 58 180 62
rect -21 -61 44 -57
rect -21 -62 -17 -61
rect 48 -67 52 58
rect 144 49 148 53
rect -11 -71 52 -67
rect 56 -76 60 49
rect 164 40 168 44
rect -1 -80 60 -76
rect 64 -85 68 40
rect 112 25 116 29
rect 9 -89 68 -85
rect 72 -92 76 20
rect 112 0 116 20
rect 122 10 126 29
rect 132 25 136 29
rect 122 6 136 10
rect 132 0 136 6
rect 112 -4 122 0
rect 142 0 146 29
rect 152 25 156 29
rect 162 17 166 29
rect 152 13 166 17
rect 152 0 156 13
rect -33 -112 -29 -100
rect -13 -105 -9 -100
rect -33 -123 -29 -117
rect -23 -109 -9 -105
rect -23 -123 -19 -109
rect -13 -123 -9 -117
rect -3 -123 1 -100
rect 21 -100 26 -96
rect 47 -96 76 -92
rect 90 -19 138 -15
rect 31 -100 41 -96
rect 7 -105 11 -100
rect 7 -109 21 -105
rect 7 -123 11 -117
rect 17 -123 21 -109
rect 27 -123 31 -117
rect 37 -114 41 -100
rect 47 -102 51 -96
rect 57 -114 61 -110
rect 90 -111 94 -19
rect 98 -28 148 -24
rect 37 -118 49 -114
rect 57 -118 78 -114
rect 37 -123 41 -118
rect 57 -123 61 -118
rect 98 -120 102 -28
rect 106 -37 158 -33
rect -35 -134 -31 -130
rect 47 -131 51 -127
rect 106 -130 110 -37
rect 162 -38 166 -8
rect 120 -46 124 -42
rect 176 -48 180 58
rect 134 -52 180 -48
rect 243 49 284 53
rect 134 -53 138 -52
rect 184 -58 188 49
rect 263 40 267 44
rect 144 -62 188 -58
rect 192 -67 196 40
rect 231 25 235 29
rect 154 -71 196 -67
rect 200 -76 204 20
rect 231 7 235 20
rect 241 17 245 29
rect 251 25 255 29
rect 241 13 255 17
rect 251 7 255 13
rect 231 3 241 7
rect 261 7 265 29
rect 122 -94 126 -82
rect 142 -87 146 -82
rect 122 -105 126 -99
rect 132 -91 146 -87
rect 166 -82 169 -78
rect 174 -82 176 -78
rect 132 -105 136 -91
rect 142 -105 146 -99
rect 152 -105 156 -82
rect 162 -105 166 -99
rect 172 -96 176 -82
rect 182 -79 204 -76
rect 217 -12 257 -8
rect 182 -84 186 -79
rect 217 -87 221 -12
rect 225 -21 267 -17
rect 192 -96 196 -92
rect 172 -100 184 -96
rect 192 -100 205 -96
rect 225 -97 229 -21
rect 271 -25 275 -1
rect 239 -30 243 -26
rect 280 -33 284 49
rect 344 42 366 46
rect 253 -37 284 -33
rect 253 -38 257 -37
rect 288 -43 292 40
rect 332 25 336 31
rect 263 -47 292 -43
rect 296 -52 300 20
rect 332 13 336 20
rect 342 13 346 31
rect 241 -70 245 -58
rect 261 -63 265 -58
rect 241 -81 245 -75
rect 251 -67 265 -63
rect 275 -58 278 -54
rect 251 -81 255 -67
rect 261 -81 265 -75
rect 271 -72 275 -58
rect 287 -55 300 -52
rect 316 -6 348 -2
rect 352 -4 356 5
rect 287 -60 291 -55
rect 316 -61 320 -6
rect 330 -15 334 -11
rect 362 -19 366 42
rect 344 -23 366 -19
rect 344 -24 348 -23
rect 370 -26 374 21
rect 368 -29 374 -26
rect 356 -35 359 -31
rect 332 -43 336 -35
rect 352 -40 356 -35
rect 332 -54 336 -48
rect 342 -43 356 -40
rect 368 -36 372 -29
rect 342 -54 346 -43
rect 359 -48 363 -36
rect 378 -48 382 -44
rect 359 -52 370 -48
rect 378 -52 388 -48
rect 378 -56 382 -52
rect 365 -60 368 -56
rect 316 -65 334 -61
rect 297 -72 301 -68
rect 271 -76 289 -72
rect 297 -76 308 -72
rect 271 -81 275 -76
rect 297 -81 301 -76
rect 239 -92 243 -88
rect 287 -89 291 -85
rect 172 -105 176 -100
rect 192 -105 196 -100
rect 225 -101 263 -97
rect 120 -116 124 -112
rect 182 -113 186 -109
rect 140 -125 144 -121
rect 106 -134 164 -130
rect -15 -143 -11 -139
rect 5 -152 9 -148
rect -49 -161 29 -157
<< m2contact >>
rect -7 58 -2 63
rect 13 49 18 54
rect 32 40 37 45
rect -44 20 -39 25
rect -24 20 -19 25
rect -4 20 1 25
rect 16 20 21 25
rect -73 -134 -68 -129
rect -65 -143 -60 -138
rect -57 -152 -52 -147
rect 17 -54 22 -49
rect 47 58 52 63
rect 55 49 60 54
rect 148 49 153 54
rect 63 40 68 45
rect 168 40 173 45
rect 71 20 76 25
rect 111 20 116 25
rect 131 20 136 25
rect 151 20 156 25
rect -34 -117 -29 -112
rect -14 -117 -9 -112
rect 26 -100 31 -95
rect 6 -117 11 -112
rect 26 -117 31 -112
rect 90 -116 95 -111
rect 98 -125 103 -120
rect -40 -135 -35 -130
rect 46 -136 51 -131
rect 162 -43 167 -38
rect 184 49 189 54
rect 191 40 196 45
rect 267 40 272 45
rect 199 20 204 25
rect 230 20 235 25
rect 250 20 255 25
rect 121 -99 126 -94
rect 169 -82 174 -77
rect 141 -99 146 -94
rect 161 -99 166 -94
rect 217 -92 222 -87
rect 271 -30 276 -25
rect 287 40 292 45
rect 295 20 300 25
rect 332 20 337 25
rect 240 -75 245 -70
rect 260 -75 265 -70
rect 278 -59 283 -54
rect 352 -9 357 -4
rect 369 21 374 26
rect 331 -48 336 -43
rect 359 -36 364 -31
rect 360 -60 365 -55
rect 234 -93 239 -88
rect 286 -94 291 -89
rect 115 -117 120 -112
rect 181 -118 186 -113
rect 135 -126 140 -121
rect -20 -144 -15 -139
rect 0 -153 5 -148
<< metal2 >>
rect -2 58 47 62
rect 18 49 55 53
rect 153 49 184 53
rect 37 40 63 44
rect 173 40 191 44
rect 272 40 287 44
rect -39 20 -24 24
rect -19 20 -4 24
rect 1 20 16 24
rect 21 20 71 24
rect 116 20 131 24
rect 136 20 151 24
rect 156 20 199 24
rect 235 20 250 24
rect 255 20 295 24
rect 337 21 369 25
rect 352 -25 356 -9
rect 352 -29 364 -25
rect 272 -38 276 -30
rect 359 -31 364 -29
rect 167 -43 174 -39
rect 272 -42 283 -38
rect 22 -54 31 -50
rect 27 -95 31 -54
rect 170 -77 174 -43
rect 279 -54 283 -42
rect 336 -48 351 -44
rect 347 -56 351 -48
rect 347 -60 360 -56
rect 245 -75 260 -71
rect 222 -92 234 -88
rect 256 -89 260 -75
rect 256 -93 286 -89
rect 126 -99 141 -95
rect 146 -99 161 -95
rect -29 -117 -14 -113
rect -9 -117 6 -113
rect 11 -117 26 -113
rect 95 -116 115 -112
rect 157 -113 161 -99
rect 157 -117 181 -113
rect -68 -134 -40 -130
rect 2 -131 6 -117
rect 103 -125 135 -121
rect 2 -135 46 -131
rect -60 -143 -20 -139
rect -52 -152 0 -148
<< labels >>
rlabel pdcontact -31 -7 -30 -5 1 vdd
rlabel ndcontact -31 -99 -30 -98 1 gnd
rlabel metal1 -20 -18 -18 -17 1 g0
rlabel metal1 -10 -27 -8 -26 1 g1
rlabel metal1 0 -36 2 -35 1 g2
rlabel metal1 10 -45 12 -44 1 g3
rlabel metal1 -20 -61 -18 -60 1 p0
rlabel metal1 0 -79 2 -78 1 p2
rlabel metal1 10 -88 12 -87 1 p3
rlabel metal1 -10 -70 -8 -69 1 p1
rlabel metal1 75 -116 77 -115 7 c4
rlabel metal1 38 -117 41 -116 1 c4_bar
rlabel metal1 -34 -53 -32 -52 1 c0
rlabel pdcontact -22 -6 -21 -4 1 u40
rlabel pdcontact -12 -6 -11 -4 1 u41
rlabel pdcontact -2 -6 -1 -4 1 u42
rlabel pdcontact 8 -6 9 -4 1 u43
rlabel ndcontact -22 -99 -21 -98 1 g40
rlabel ndcontact -12 -99 -11 -98 1 g41
rlabel ndcontact -2 -99 -1 -98 1 g42
rlabel ndcontact 8 -99 9 -98 1 g43
rlabel pdcontact 124 -7 125 -5 1 vdd
rlabel metal1 135 -18 137 -17 1 g0
rlabel metal1 145 -27 147 -26 1 g1
rlabel metal1 155 -36 157 -35 1 g2
rlabel metal1 121 -45 123 -44 1 c0
rlabel metal1 135 -52 137 -51 1 p0
rlabel metal1 155 -70 157 -69 1 p2
rlabel metal1 145 -61 147 -60 1 p1
rlabel ndcontact 124 -81 125 -80 1 gnd
rlabel pdcontact 133 -6 134 -4 1 u30
rlabel pdcontact 143 -6 144 -4 1 u31
rlabel pdcontact 153 -6 154 -4 1 u32
rlabel ndcontact 133 -81 134 -80 1 g30
rlabel ndcontact 143 -81 144 -80 1 g31
rlabel ndcontact 153 -81 154 -80 1 g32
rlabel metal1 176 -99 179 -98 1 c3_bar
rlabel metal1 201 -100 203 -99 1 c3
rlabel metal1 304 -76 306 -75 1 c2
rlabel metal1 277 -75 279 -74 1 c2_bar
rlabel pdcontact 262 1 263 3 1 u21
rlabel pdcontact 252 1 253 3 1 u20
rlabel ndcontact 262 -57 263 -56 1 d21
rlabel ndcontact 252 -57 253 -56 1 d20
rlabel ndcontact 243 -57 244 -56 1 gnd
rlabel metal1 264 -46 266 -45 1 p1
rlabel metal1 254 -37 256 -36 1 p0
rlabel metal1 240 -29 242 -28 1 c0
rlabel metal1 264 -20 266 -19 1 g1
rlabel metal1 254 -11 256 -10 1 g0
rlabel pdcontact 243 0 244 2 1 vdd
rlabel pdcontact 334 6 335 8 1 vdd
rlabel metal1 345 -5 347 -4 1 g0
rlabel metal1 331 -14 333 -13 1 c0
rlabel metal1 345 -23 347 -22 1 p0
rlabel ndcontact 334 -34 335 -33 1 gnd
rlabel pdcontact 343 7 344 9 1 u10
rlabel ndcontact 343 -34 344 -33 1 d10
rlabel metal1 360 -51 362 -50 1 c1_bar
rlabel metal1 386 -51 388 -50 7 c1
<< end >>

magic
tech scmos
timestamp 1619482272
<< nwell >>
rect -58 -60 -4 -40
rect 12 -49 44 -7
rect 100 -60 154 -40
rect 170 -49 202 -7
rect -58 -158 -4 -138
rect 12 -147 44 -105
rect 100 -158 154 -138
rect 170 -147 202 -105
<< ntransistor >>
rect -47 -70 -45 -66
rect -17 -70 -15 -66
rect 23 -67 25 -63
rect 31 -67 33 -63
rect 111 -70 113 -66
rect 141 -70 143 -66
rect 181 -67 183 -63
rect 189 -67 191 -63
rect 23 -89 25 -85
rect 31 -89 33 -85
rect 181 -89 183 -85
rect 189 -89 191 -85
rect -47 -168 -45 -164
rect -17 -168 -15 -164
rect 23 -165 25 -161
rect 31 -165 33 -161
rect 111 -168 113 -164
rect 141 -168 143 -164
rect 181 -165 183 -161
rect 189 -165 191 -161
rect 23 -187 25 -183
rect 31 -187 33 -183
rect 181 -187 183 -183
rect 189 -187 191 -183
<< ptransistor >>
rect 23 -21 25 -13
rect 31 -21 33 -13
rect 181 -21 183 -13
rect 189 -21 191 -13
rect 23 -43 25 -35
rect 31 -43 33 -35
rect 181 -43 183 -35
rect 189 -43 191 -35
rect -47 -54 -45 -46
rect -17 -54 -15 -46
rect 111 -54 113 -46
rect 141 -54 143 -46
rect 23 -119 25 -111
rect 31 -119 33 -111
rect 181 -119 183 -111
rect 189 -119 191 -111
rect 23 -141 25 -133
rect 31 -141 33 -133
rect 181 -141 183 -133
rect 189 -141 191 -133
rect -47 -152 -45 -144
rect -17 -152 -15 -144
rect 111 -152 113 -144
rect 141 -152 143 -144
<< ndiffusion >>
rect -48 -70 -47 -66
rect -45 -70 -44 -66
rect -18 -70 -17 -66
rect -15 -70 -14 -66
rect 22 -67 23 -63
rect 25 -67 26 -63
rect 30 -67 31 -63
rect 33 -67 34 -63
rect 110 -70 111 -66
rect 113 -70 114 -66
rect 140 -70 141 -66
rect 143 -70 144 -66
rect 180 -67 181 -63
rect 183 -67 184 -63
rect 188 -67 189 -63
rect 191 -67 192 -63
rect 22 -89 23 -85
rect 25 -89 26 -85
rect 30 -89 31 -85
rect 33 -89 34 -85
rect 180 -89 181 -85
rect 183 -89 184 -85
rect 188 -89 189 -85
rect 191 -89 192 -85
rect -48 -168 -47 -164
rect -45 -168 -44 -164
rect -18 -168 -17 -164
rect -15 -168 -14 -164
rect 22 -165 23 -161
rect 25 -165 26 -161
rect 30 -165 31 -161
rect 33 -165 34 -161
rect 110 -168 111 -164
rect 113 -168 114 -164
rect 140 -168 141 -164
rect 143 -168 144 -164
rect 180 -165 181 -161
rect 183 -165 184 -161
rect 188 -165 189 -161
rect 191 -165 192 -161
rect 22 -187 23 -183
rect 25 -187 26 -183
rect 30 -187 31 -183
rect 33 -187 34 -183
rect 180 -187 181 -183
rect 183 -187 184 -183
rect 188 -187 189 -183
rect 191 -187 192 -183
<< pdiffusion >>
rect 22 -21 23 -13
rect 25 -21 26 -13
rect 30 -21 31 -13
rect 33 -21 34 -13
rect 180 -21 181 -13
rect 183 -21 184 -13
rect 188 -21 189 -13
rect 191 -21 192 -13
rect 22 -43 23 -35
rect 25 -43 26 -35
rect 30 -43 31 -35
rect 33 -43 34 -35
rect 180 -43 181 -35
rect 183 -43 184 -35
rect 188 -43 189 -35
rect 191 -43 192 -35
rect -48 -54 -47 -46
rect -45 -54 -44 -46
rect -18 -54 -17 -46
rect -15 -54 -14 -46
rect 110 -54 111 -46
rect 113 -54 114 -46
rect 140 -54 141 -46
rect 143 -54 144 -46
rect 22 -119 23 -111
rect 25 -119 26 -111
rect 30 -119 31 -111
rect 33 -119 34 -111
rect 180 -119 181 -111
rect 183 -119 184 -111
rect 188 -119 189 -111
rect 191 -119 192 -111
rect 22 -141 23 -133
rect 25 -141 26 -133
rect 30 -141 31 -133
rect 33 -141 34 -133
rect 180 -141 181 -133
rect 183 -141 184 -133
rect 188 -141 189 -133
rect 191 -141 192 -133
rect -48 -152 -47 -144
rect -45 -152 -44 -144
rect -18 -152 -17 -144
rect -15 -152 -14 -144
rect 110 -152 111 -144
rect 113 -152 114 -144
rect 140 -152 141 -144
rect 143 -152 144 -144
<< ndcontact >>
rect -52 -70 -48 -66
rect -44 -70 -40 -66
rect -22 -70 -18 -66
rect -14 -70 -10 -66
rect 18 -67 22 -63
rect 26 -67 30 -63
rect 34 -67 38 -63
rect 106 -70 110 -66
rect 114 -70 118 -66
rect 136 -70 140 -66
rect 144 -70 148 -66
rect 176 -67 180 -63
rect 184 -67 188 -63
rect 192 -67 196 -63
rect 18 -89 22 -85
rect 26 -89 30 -85
rect 34 -89 38 -85
rect 176 -89 180 -85
rect 184 -89 188 -85
rect 192 -89 196 -85
rect -52 -168 -48 -164
rect -44 -168 -40 -164
rect -22 -168 -18 -164
rect -14 -168 -10 -164
rect 18 -165 22 -161
rect 26 -165 30 -161
rect 34 -165 38 -161
rect 106 -168 110 -164
rect 114 -168 118 -164
rect 136 -168 140 -164
rect 144 -168 148 -164
rect 176 -165 180 -161
rect 184 -165 188 -161
rect 192 -165 196 -161
rect 18 -187 22 -183
rect 26 -187 30 -183
rect 34 -187 38 -183
rect 176 -187 180 -183
rect 184 -187 188 -183
rect 192 -187 196 -183
<< pdcontact >>
rect 18 -21 22 -13
rect 26 -21 30 -13
rect 34 -21 38 -13
rect 176 -21 180 -13
rect 184 -21 188 -13
rect 192 -21 196 -13
rect 18 -43 22 -35
rect 26 -43 30 -35
rect 34 -43 38 -35
rect 176 -43 180 -35
rect 184 -43 188 -35
rect 192 -43 196 -35
rect -52 -54 -48 -46
rect -44 -54 -40 -46
rect -22 -54 -18 -46
rect -14 -54 -10 -46
rect 106 -54 110 -46
rect 114 -54 118 -46
rect 136 -54 140 -46
rect 144 -54 148 -46
rect 18 -119 22 -111
rect 26 -119 30 -111
rect 34 -119 38 -111
rect 176 -119 180 -111
rect 184 -119 188 -111
rect 192 -119 196 -111
rect 18 -141 22 -133
rect 26 -141 30 -133
rect 34 -141 38 -133
rect 176 -141 180 -133
rect 184 -141 188 -133
rect 192 -141 196 -133
rect -52 -152 -48 -144
rect -44 -152 -40 -144
rect -22 -152 -18 -144
rect -14 -152 -10 -144
rect 106 -152 110 -144
rect 114 -152 118 -144
rect 136 -152 140 -144
rect 144 -152 148 -144
<< polysilicon >>
rect 23 -13 25 -10
rect 31 -13 33 -10
rect 181 -13 183 -10
rect 189 -13 191 -10
rect 23 -28 25 -21
rect 31 -28 33 -21
rect 181 -28 183 -21
rect 189 -28 191 -21
rect 23 -35 25 -32
rect 31 -35 33 -32
rect 181 -35 183 -32
rect 189 -35 191 -32
rect -47 -46 -45 -43
rect -17 -46 -15 -43
rect -47 -66 -45 -54
rect -17 -66 -15 -54
rect 23 -63 25 -43
rect 31 -51 33 -43
rect 111 -46 113 -43
rect 141 -46 143 -43
rect 31 -63 33 -55
rect 111 -66 113 -54
rect 141 -66 143 -54
rect 181 -63 183 -43
rect 189 -51 191 -43
rect 189 -63 191 -55
rect 23 -70 25 -67
rect 31 -70 33 -67
rect 181 -70 183 -67
rect 189 -70 191 -67
rect -47 -73 -45 -70
rect -17 -73 -15 -70
rect 111 -73 113 -70
rect 141 -73 143 -70
rect 23 -85 25 -78
rect 31 -85 33 -78
rect 181 -85 183 -78
rect 189 -85 191 -78
rect 23 -92 25 -89
rect 31 -92 33 -89
rect 181 -92 183 -89
rect 189 -92 191 -89
rect 23 -111 25 -108
rect 31 -111 33 -108
rect 181 -111 183 -108
rect 189 -111 191 -108
rect 23 -126 25 -119
rect 31 -126 33 -119
rect 181 -126 183 -119
rect 189 -126 191 -119
rect 23 -133 25 -130
rect 31 -133 33 -130
rect 181 -133 183 -130
rect 189 -133 191 -130
rect -47 -144 -45 -141
rect -17 -144 -15 -141
rect -47 -164 -45 -152
rect -17 -164 -15 -152
rect 23 -161 25 -141
rect 31 -149 33 -141
rect 111 -144 113 -141
rect 141 -144 143 -141
rect 31 -161 33 -153
rect 111 -164 113 -152
rect 141 -164 143 -152
rect 181 -161 183 -141
rect 189 -149 191 -141
rect 189 -161 191 -153
rect 23 -168 25 -165
rect 31 -168 33 -165
rect 181 -168 183 -165
rect 189 -168 191 -165
rect -47 -171 -45 -168
rect -17 -171 -15 -168
rect 111 -171 113 -168
rect 141 -171 143 -168
rect 23 -183 25 -176
rect 31 -183 33 -176
rect 181 -183 183 -176
rect 189 -183 191 -176
rect 23 -190 25 -187
rect 31 -190 33 -187
rect 181 -190 183 -187
rect 189 -190 191 -187
<< polycontact >>
rect 19 -28 23 -24
rect 33 -28 37 -24
rect 177 -28 181 -24
rect 191 -28 195 -24
rect -51 -62 -47 -58
rect -21 -62 -17 -58
rect 19 -57 23 -53
rect 33 -50 37 -46
rect 33 -60 37 -56
rect 107 -62 111 -58
rect 137 -62 141 -58
rect 177 -57 181 -53
rect 191 -50 195 -46
rect 191 -60 195 -56
rect 19 -82 23 -78
rect 33 -82 37 -78
rect 177 -82 181 -78
rect 191 -82 195 -78
rect 19 -126 23 -122
rect 33 -126 37 -122
rect 177 -126 181 -122
rect 191 -126 195 -122
rect -51 -160 -47 -156
rect -21 -160 -17 -156
rect 19 -155 23 -151
rect 33 -148 37 -144
rect 33 -158 37 -154
rect 107 -160 111 -156
rect 137 -160 141 -156
rect 177 -155 181 -151
rect 191 -148 195 -144
rect 191 -158 195 -154
rect 19 -180 23 -176
rect 33 -180 37 -176
rect 177 -180 181 -176
rect 191 -180 195 -176
<< metal1 >>
rect -91 38 -45 42
rect -91 29 -52 33
rect -91 20 -64 24
rect -91 11 -82 15
rect -56 15 -52 29
rect -49 24 -45 38
rect 227 37 247 41
rect 236 28 247 32
rect -49 20 94 24
rect 115 20 247 24
rect -56 11 76 15
rect 123 11 247 15
rect -91 3 247 6
rect -77 -111 -73 3
rect -57 -39 -53 3
rect 0 -35 4 3
rect 18 -13 22 3
rect 57 -15 61 -1
rect 38 -19 61 -15
rect 16 -28 19 -24
rect 37 -28 40 -24
rect 0 -39 18 -35
rect -57 -42 -18 -39
rect -69 -49 -64 -45
rect -52 -46 -48 -42
rect -22 -46 -18 -42
rect 57 -37 61 -19
rect 38 -41 61 -37
rect 37 -50 40 -46
rect -44 -57 -40 -54
rect -69 -62 -60 -58
rect -55 -62 -51 -58
rect -44 -66 -40 -62
rect -24 -62 -21 -58
rect -14 -66 -10 -54
rect 15 -57 19 -53
rect 37 -60 40 -56
rect 57 -63 61 -41
rect 0 -67 18 -63
rect 38 -67 61 -63
rect -52 -85 -48 -70
rect -22 -85 -18 -70
rect 0 -85 4 -67
rect 19 -78 23 -76
rect 33 -78 37 -76
rect 57 -85 61 -67
rect -70 -88 18 -85
rect -65 -89 18 -88
rect 38 -89 61 -85
rect 81 -111 85 3
rect 101 -39 105 3
rect 158 -35 162 3
rect 176 -13 180 3
rect 196 -19 219 -15
rect 174 -28 177 -24
rect 195 -28 198 -24
rect 158 -39 176 -35
rect 101 -42 140 -39
rect 89 -49 94 -45
rect 106 -46 110 -42
rect 136 -46 140 -42
rect 215 -37 219 -19
rect 196 -41 219 -37
rect 195 -50 198 -46
rect 215 -51 219 -41
rect 222 -51 226 -8
rect 114 -57 118 -54
rect 89 -62 98 -58
rect 103 -62 107 -58
rect 114 -66 118 -62
rect 134 -62 137 -58
rect 144 -66 148 -54
rect 173 -57 177 -53
rect 215 -55 226 -51
rect 195 -60 198 -56
rect 215 -63 219 -55
rect 158 -67 176 -63
rect 196 -67 219 -63
rect 106 -85 110 -70
rect 136 -85 140 -70
rect 158 -85 162 -67
rect 177 -78 181 -76
rect 191 -78 195 -76
rect 215 -85 219 -67
rect 88 -88 176 -85
rect 93 -89 176 -88
rect 196 -89 219 -85
rect -77 -115 18 -111
rect -57 -137 -53 -115
rect 0 -133 4 -115
rect 38 -117 61 -113
rect 81 -115 176 -111
rect 16 -126 19 -122
rect 37 -126 40 -122
rect 0 -137 18 -133
rect -57 -140 -18 -137
rect -69 -147 -64 -143
rect -52 -144 -48 -140
rect -22 -144 -18 -140
rect 57 -135 61 -117
rect 38 -139 61 -135
rect 37 -148 40 -144
rect 57 -148 61 -139
rect 101 -137 105 -115
rect 158 -133 162 -115
rect 196 -117 219 -113
rect 174 -126 177 -122
rect 195 -126 198 -122
rect 158 -137 176 -133
rect 101 -140 140 -137
rect 89 -147 94 -143
rect 106 -144 110 -140
rect 136 -144 140 -140
rect 215 -135 219 -117
rect 196 -139 219 -135
rect -44 -155 -40 -152
rect -69 -160 -60 -156
rect -55 -160 -51 -156
rect -44 -164 -40 -160
rect -24 -160 -21 -156
rect -14 -164 -10 -152
rect 15 -155 19 -151
rect 57 -153 62 -148
rect 195 -148 198 -144
rect 215 -149 219 -139
rect 232 -149 236 -8
rect 37 -158 40 -154
rect 57 -161 61 -153
rect 114 -155 118 -152
rect 89 -160 98 -156
rect 103 -160 107 -156
rect 0 -165 18 -161
rect 38 -165 61 -161
rect 114 -164 118 -160
rect 134 -160 137 -156
rect 144 -164 148 -152
rect 173 -155 177 -151
rect 215 -153 236 -149
rect 195 -158 198 -154
rect 215 -161 219 -153
rect -91 -205 -74 -202
rect -52 -202 -48 -168
rect -22 -202 -18 -168
rect 0 -202 4 -165
rect 19 -176 23 -174
rect 33 -176 37 -174
rect 57 -183 61 -165
rect 38 -187 61 -183
rect 158 -165 176 -161
rect 196 -165 219 -161
rect 18 -202 22 -187
rect -69 -205 84 -202
rect 106 -202 110 -168
rect 136 -202 140 -168
rect 158 -202 162 -165
rect 177 -176 181 -174
rect 191 -176 195 -174
rect 215 -183 219 -165
rect 196 -187 219 -183
rect 176 -202 180 -187
rect 89 -205 247 -202
rect -91 -214 -59 -210
rect -51 -214 99 -210
rect -91 -223 -85 -219
rect -51 -228 -46 -214
rect -91 -232 -46 -228
rect -42 -223 71 -219
rect -42 -237 -38 -223
rect -91 -241 -38 -237
<< m2contact >>
rect 222 36 227 41
rect 231 28 236 33
rect 110 20 115 25
rect 118 10 123 15
rect 61 -5 66 0
rect 40 -51 45 -46
rect -60 -63 -55 -58
rect 10 -57 15 -52
rect -10 -63 -5 -58
rect 33 -76 38 -71
rect -70 -93 -65 -88
rect 222 -8 227 -3
rect 231 -8 236 -3
rect 198 -51 203 -46
rect 98 -63 103 -58
rect 168 -57 173 -52
rect 148 -63 153 -58
rect 191 -76 196 -71
rect 88 -93 93 -88
rect 40 -149 45 -144
rect -60 -161 -55 -156
rect 10 -155 15 -150
rect 62 -153 67 -148
rect 198 -149 203 -144
rect -10 -161 -5 -156
rect 98 -161 103 -156
rect 168 -155 173 -150
rect 148 -161 153 -156
rect -74 -205 -69 -200
rect 33 -174 38 -169
rect 84 -205 89 -200
rect 191 -174 196 -169
rect -59 -214 -54 -209
rect 99 -214 104 -209
rect -85 -223 -80 -218
rect 71 -223 76 -218
<< metal2 >>
rect -5 -7 56 -3
rect 110 -1 114 20
rect 66 -5 114 -1
rect -5 -63 -1 -7
rect 52 -46 56 -7
rect 118 -9 122 10
rect 222 -3 226 36
rect 232 -3 236 28
rect 45 -50 56 -46
rect -59 -79 -55 -63
rect 10 -79 14 -57
rect 52 -72 56 -50
rect 38 -76 56 -72
rect 63 -13 122 -9
rect 153 -7 214 -3
rect -87 -83 14 -79
rect -87 -111 -83 -83
rect -87 -114 -81 -111
rect -85 -218 -81 -114
rect -70 -119 -66 -93
rect -77 -123 -66 -119
rect -5 -105 56 -101
rect -77 -197 -73 -123
rect -5 -161 -1 -105
rect 52 -144 56 -105
rect 45 -148 56 -144
rect 63 -148 67 -13
rect 153 -63 157 -7
rect 210 -46 214 -7
rect 203 -50 214 -46
rect 99 -79 103 -63
rect 168 -79 172 -57
rect 210 -72 214 -50
rect 196 -76 214 -72
rect -59 -183 -55 -161
rect 10 -183 14 -155
rect 52 -170 56 -148
rect 71 -83 172 -79
rect 38 -174 56 -170
rect -59 -187 14 -183
rect -77 -200 -69 -197
rect -59 -209 -55 -187
rect 71 -218 75 -83
rect 88 -119 92 -93
rect 81 -123 92 -119
rect 153 -105 214 -101
rect 81 -190 85 -123
rect 153 -161 157 -105
rect 210 -144 214 -105
rect 203 -148 214 -144
rect 99 -183 103 -161
rect 168 -183 172 -155
rect 210 -170 214 -148
rect 196 -174 214 -170
rect 99 -187 172 -183
rect 81 -194 88 -190
rect 84 -200 88 -194
rect 99 -209 103 -187
<< m123contact >>
rect -64 20 -59 25
rect 94 20 99 25
rect -82 11 -77 16
rect 76 11 81 16
rect -64 -50 -59 -45
rect -44 -62 -39 -57
rect -29 -63 -24 -58
rect 11 -29 16 -24
rect 40 -29 45 -24
rect 40 -60 45 -55
rect 18 -76 23 -71
rect -64 -148 -59 -143
rect -44 -160 -39 -155
rect -29 -161 -24 -156
rect 11 -127 16 -122
rect 40 -127 45 -122
rect 94 -50 99 -45
rect 114 -62 119 -57
rect 129 -63 134 -58
rect 169 -29 174 -24
rect 198 -29 203 -24
rect 198 -60 203 -55
rect 176 -76 181 -71
rect 40 -158 45 -153
rect 18 -174 23 -169
rect 94 -148 99 -143
rect 114 -160 119 -155
rect 129 -161 134 -156
rect 169 -127 174 -122
rect 198 -127 203 -122
rect 198 -158 203 -153
rect 176 -174 181 -169
<< metal3 >>
rect -82 -105 -78 11
rect -64 -45 -60 20
rect -37 -29 11 -24
rect 45 -29 51 -25
rect -64 -93 -61 -50
rect -37 -57 -33 -29
rect -39 -61 -33 -57
rect -29 -93 -25 -63
rect 5 -71 9 -29
rect 47 -55 51 -29
rect 45 -60 51 -55
rect 5 -76 18 -71
rect 41 -93 45 -60
rect -64 -97 45 -93
rect 76 -105 80 11
rect 94 -45 98 20
rect 121 -29 169 -24
rect 203 -29 209 -25
rect 94 -93 97 -50
rect 121 -57 125 -29
rect 119 -61 125 -57
rect 129 -93 133 -63
rect 163 -71 167 -29
rect 205 -55 209 -29
rect 203 -60 209 -55
rect 163 -76 176 -71
rect 199 -93 203 -60
rect 94 -97 203 -93
rect -82 -109 -60 -105
rect 76 -109 98 -105
rect -64 -143 -60 -109
rect -37 -127 11 -122
rect 45 -127 51 -123
rect -64 -193 -61 -148
rect -37 -155 -33 -127
rect -39 -159 -33 -155
rect -29 -193 -25 -161
rect 5 -169 9 -127
rect 47 -153 51 -127
rect 45 -158 51 -153
rect 94 -143 98 -109
rect 121 -127 169 -122
rect 203 -127 209 -123
rect 5 -174 18 -169
rect 41 -193 45 -158
rect -64 -197 45 -193
rect 94 -193 97 -148
rect 121 -155 125 -127
rect 119 -159 125 -155
rect 129 -193 133 -161
rect 163 -169 167 -127
rect 205 -153 209 -127
rect 203 -158 209 -153
rect 163 -174 176 -169
rect 199 -193 203 -158
rect 94 -197 203 -193
<< labels >>
rlabel metal1 1 -204 3 -203 1 gnd
rlabel metal1 -90 -204 -88 -203 3 gnd
rlabel metal1 236 -205 238 -204 1 gnd
rlabel metal1 159 -204 161 -203 1 gnd
rlabel metal1 159 4 161 5 5 vdd
rlabel metal1 240 3 242 4 1 vdd
rlabel metal1 -89 4 -87 5 3 vdd
rlabel metal1 1 4 3 5 5 vdd
rlabel pdcontact 27 -118 28 -116 1 xs00
rlabel pdcontact 27 -140 28 -138 1 xs01
rlabel ndcontact 27 -164 28 -163 1 xs02
rlabel ndcontact 27 -186 28 -185 1 xs03
rlabel metal1 -89 12 -87 13 3 p0
rlabel metal1 -89 21 -87 22 3 p1
rlabel metal1 -89 30 -87 31 3 p2
rlabel metal1 -89 40 -87 41 4 p3
rlabel metal1 -90 -213 -88 -212 3 c0
rlabel metal1 -90 -222 -88 -221 3 c1
rlabel metal1 -90 -231 -88 -230 3 c2
rlabel metal1 -90 -240 -88 -239 2 c3
rlabel metal1 -43 -163 -41 -162 1 c0_bar
rlabel metal1 -13 -163 -11 -162 1 p0_bar
rlabel metal1 -43 -65 -41 -64 1 c1_bar
rlabel metal1 -13 -65 -11 -64 1 p1_bar
rlabel metal1 115 -163 117 -162 1 c2_bar
rlabel metal1 145 -163 147 -162 1 p2_bar
rlabel metal1 115 -65 117 -64 1 c3_bar
rlabel metal1 145 -65 147 -64 1 p3_bar
rlabel pdcontact 27 -20 28 -18 1 xs10
rlabel pdcontact 27 -42 28 -40 1 xs11
rlabel ndcontact 27 -66 28 -65 1 xs12
rlabel ndcontact 27 -88 28 -87 1 xs13
rlabel pdcontact 185 -117 186 -116 1 xs20
rlabel pdcontact 185 -139 186 -138 1 xs21
rlabel ndcontact 185 -164 186 -163 1 xs22
rlabel ndcontact 185 -186 186 -185 1 xs23
rlabel pdcontact 185 -19 186 -18 1 xs30
rlabel pdcontact 185 -41 186 -40 1 xs31
rlabel ndcontact 185 -66 186 -65 1 xs32
rlabel ndcontact 185 -88 186 -87 1 xs33
rlabel metal1 240 12 242 13 1 s0
rlabel metal1 240 21 242 22 1 s1
rlabel metal1 240 29 242 30 1 s2
rlabel metal1 240 39 242 40 5 s3
<< end >>

magic
tech scmos
timestamp 1619564990
<< nwell >>
rect 1960 193 1984 214
rect 1991 187 2023 215
rect 2033 178 2057 198
rect 2069 187 2101 215
rect 2137 187 2169 215
rect 2179 178 2203 198
rect 2215 187 2247 215
rect -67 81 -43 102
rect -35 90 -3 118
rect 7 81 31 101
rect 43 90 75 118
rect 111 90 143 118
rect 153 81 177 101
rect 189 90 221 118
rect 233 81 257 102
rect 263 90 295 118
rect 305 81 329 101
rect 341 90 373 118
rect 409 90 441 118
rect 451 81 475 101
rect 487 90 519 118
rect 531 81 555 102
rect 561 90 593 118
rect 603 81 627 101
rect 639 90 671 118
rect 707 90 739 118
rect 749 81 773 101
rect 785 90 817 118
rect 829 81 853 102
rect 859 90 891 118
rect 901 81 925 101
rect 937 90 969 118
rect 1005 90 1037 118
rect 1047 81 1071 101
rect 1083 90 1115 118
rect 1966 81 1990 102
rect 1998 90 2030 118
rect 2040 81 2064 101
rect 2076 90 2108 118
rect 2144 90 2176 118
rect 2186 81 2210 101
rect 2222 90 2254 118
rect 2266 81 2290 102
rect 2296 90 2328 118
rect 2338 81 2362 101
rect 2374 90 2406 118
rect 2442 90 2474 118
rect 2484 81 2508 101
rect 2520 90 2552 118
rect -67 -20 -43 1
rect -35 -11 -3 17
rect 43 -11 75 17
rect 111 -11 143 17
rect 153 -20 177 0
rect 189 -11 221 17
rect 232 -5 256 16
rect 263 -11 295 17
rect 305 -20 329 0
rect 341 -11 373 17
rect 409 -11 441 17
rect 451 -20 475 0
rect 487 -11 519 17
rect 530 -5 554 16
rect 561 -11 593 17
rect 603 -20 627 0
rect 639 -11 671 17
rect 707 -11 739 17
rect 749 -20 773 0
rect 785 -11 817 17
rect 828 -5 852 16
rect 859 -11 891 17
rect 901 -20 925 0
rect 937 -11 969 17
rect 1005 -11 1037 17
rect 1047 -20 1071 0
rect 1083 -11 1115 17
rect 1966 -20 1990 1
rect 1998 -11 2030 17
rect 2040 -20 2064 0
rect 2076 -11 2108 17
rect 2144 -11 2176 17
rect 2186 -20 2210 0
rect 2222 -11 2254 17
rect 2265 -5 2289 16
rect 2296 -11 2328 17
rect 2338 -20 2362 0
rect 2374 -11 2406 17
rect 2442 -11 2474 17
rect 2484 -20 2508 0
rect 2520 -11 2552 17
<< ntransistor >>
rect 1971 183 1973 187
rect 2044 168 2046 172
rect 2190 168 2192 172
rect 2002 154 2004 162
rect 2010 154 2012 162
rect 2080 154 2082 162
rect 2088 154 2090 162
rect 2148 154 2150 162
rect 2156 154 2158 162
rect 2226 154 2228 162
rect 2234 154 2236 162
rect -56 71 -54 75
rect 18 71 20 75
rect 164 71 166 75
rect 244 71 246 75
rect 316 71 318 75
rect 462 71 464 75
rect 542 71 544 75
rect 614 71 616 75
rect 760 71 762 75
rect 840 71 842 75
rect 912 71 914 75
rect 1058 71 1060 75
rect 1977 71 1979 75
rect 2051 71 2053 75
rect 2197 71 2199 75
rect 2277 71 2279 75
rect 2349 71 2351 75
rect 2495 71 2497 75
rect -24 57 -22 65
rect -16 57 -14 65
rect 54 57 56 65
rect 62 57 64 65
rect 122 57 124 65
rect 130 57 132 65
rect 200 57 202 65
rect 208 57 210 65
rect 274 57 276 65
rect 282 57 284 65
rect 352 57 354 65
rect 360 57 362 65
rect 420 57 422 65
rect 428 57 430 65
rect 498 57 500 65
rect 506 57 508 65
rect 572 57 574 65
rect 580 57 582 65
rect 650 57 652 65
rect 658 57 660 65
rect 718 57 720 65
rect 726 57 728 65
rect 796 57 798 65
rect 804 57 806 65
rect 870 57 872 65
rect 878 57 880 65
rect 948 57 950 65
rect 956 57 958 65
rect 1016 57 1018 65
rect 1024 57 1026 65
rect 1094 57 1096 65
rect 1102 57 1104 65
rect 2009 57 2011 65
rect 2017 57 2019 65
rect 2087 57 2089 65
rect 2095 57 2097 65
rect 2155 57 2157 65
rect 2163 57 2165 65
rect 2233 57 2235 65
rect 2241 57 2243 65
rect 2307 57 2309 65
rect 2315 57 2317 65
rect 2385 57 2387 65
rect 2393 57 2395 65
rect 2453 57 2455 65
rect 2461 57 2463 65
rect 2531 57 2533 65
rect 2539 57 2541 65
rect -56 -30 -54 -26
rect 18 -30 20 -26
rect 164 -30 166 -26
rect 243 -15 245 -11
rect 316 -30 318 -26
rect 462 -30 464 -26
rect 541 -15 543 -11
rect 614 -30 616 -26
rect 760 -30 762 -26
rect 839 -15 841 -11
rect 912 -30 914 -26
rect 1058 -30 1060 -26
rect 1977 -30 1979 -26
rect 2051 -30 2053 -26
rect 2197 -30 2199 -26
rect 2276 -15 2278 -11
rect 2349 -30 2351 -26
rect 2495 -30 2497 -26
rect -24 -44 -22 -36
rect -16 -44 -14 -36
rect 54 -44 56 -36
rect 62 -44 64 -36
rect 122 -44 124 -36
rect 130 -44 132 -36
rect 200 -44 202 -36
rect 208 -44 210 -36
rect 274 -44 276 -36
rect 282 -44 284 -36
rect 352 -44 354 -36
rect 360 -44 362 -36
rect 420 -44 422 -36
rect 428 -44 430 -36
rect 498 -44 500 -36
rect 506 -44 508 -36
rect 572 -44 574 -36
rect 580 -44 582 -36
rect 650 -44 652 -36
rect 658 -44 660 -36
rect 718 -44 720 -36
rect 726 -44 728 -36
rect 796 -44 798 -36
rect 804 -44 806 -36
rect 870 -44 872 -36
rect 878 -44 880 -36
rect 948 -44 950 -36
rect 956 -44 958 -36
rect 1016 -44 1018 -36
rect 1024 -44 1026 -36
rect 1094 -44 1096 -36
rect 1102 -44 1104 -36
rect 2009 -44 2011 -36
rect 2017 -44 2019 -36
rect 2087 -44 2089 -36
rect 2095 -44 2097 -36
rect 2155 -44 2157 -36
rect 2163 -44 2165 -36
rect 2233 -44 2235 -36
rect 2241 -44 2243 -36
rect 2307 -44 2309 -36
rect 2315 -44 2317 -36
rect 2385 -44 2387 -36
rect 2393 -44 2395 -36
rect 2453 -44 2455 -36
rect 2461 -44 2463 -36
rect 2531 -44 2533 -36
rect 2539 -44 2541 -36
<< ptransistor >>
rect 1971 199 1973 207
rect 2002 193 2004 209
rect 2010 193 2012 209
rect 2080 193 2082 209
rect 2088 193 2090 209
rect 2148 193 2150 209
rect 2156 193 2158 209
rect 2044 184 2046 192
rect 2226 193 2228 209
rect 2234 193 2236 209
rect 2190 184 2192 192
rect -24 96 -22 112
rect -16 96 -14 112
rect -56 87 -54 95
rect 54 96 56 112
rect 62 96 64 112
rect 122 96 124 112
rect 130 96 132 112
rect 18 87 20 95
rect 200 96 202 112
rect 208 96 210 112
rect 164 87 166 95
rect 274 96 276 112
rect 282 96 284 112
rect 244 87 246 95
rect 352 96 354 112
rect 360 96 362 112
rect 420 96 422 112
rect 428 96 430 112
rect 316 87 318 95
rect 498 96 500 112
rect 506 96 508 112
rect 462 87 464 95
rect 572 96 574 112
rect 580 96 582 112
rect 542 87 544 95
rect 650 96 652 112
rect 658 96 660 112
rect 718 96 720 112
rect 726 96 728 112
rect 614 87 616 95
rect 796 96 798 112
rect 804 96 806 112
rect 760 87 762 95
rect 870 96 872 112
rect 878 96 880 112
rect 840 87 842 95
rect 948 96 950 112
rect 956 96 958 112
rect 1016 96 1018 112
rect 1024 96 1026 112
rect 912 87 914 95
rect 1094 96 1096 112
rect 1102 96 1104 112
rect 1058 87 1060 95
rect 2009 96 2011 112
rect 2017 96 2019 112
rect 1977 87 1979 95
rect 2087 96 2089 112
rect 2095 96 2097 112
rect 2155 96 2157 112
rect 2163 96 2165 112
rect 2051 87 2053 95
rect 2233 96 2235 112
rect 2241 96 2243 112
rect 2197 87 2199 95
rect 2307 96 2309 112
rect 2315 96 2317 112
rect 2277 87 2279 95
rect 2385 96 2387 112
rect 2393 96 2395 112
rect 2453 96 2455 112
rect 2461 96 2463 112
rect 2349 87 2351 95
rect 2531 96 2533 112
rect 2539 96 2541 112
rect 2495 87 2497 95
rect -24 -5 -22 11
rect -16 -5 -14 11
rect -56 -14 -54 -6
rect 54 -5 56 11
rect 62 -5 64 11
rect 122 -5 124 11
rect 130 -5 132 11
rect 18 -14 20 -6
rect 200 -5 202 11
rect 208 -5 210 11
rect 243 1 245 9
rect 164 -14 166 -6
rect 274 -5 276 11
rect 282 -5 284 11
rect 352 -5 354 11
rect 360 -5 362 11
rect 420 -5 422 11
rect 428 -5 430 11
rect 316 -14 318 -6
rect 498 -5 500 11
rect 506 -5 508 11
rect 541 1 543 9
rect 462 -14 464 -6
rect 572 -5 574 11
rect 580 -5 582 11
rect 650 -5 652 11
rect 658 -5 660 11
rect 718 -5 720 11
rect 726 -5 728 11
rect 614 -14 616 -6
rect 796 -5 798 11
rect 804 -5 806 11
rect 839 1 841 9
rect 760 -14 762 -6
rect 870 -5 872 11
rect 878 -5 880 11
rect 948 -5 950 11
rect 956 -5 958 11
rect 1016 -5 1018 11
rect 1024 -5 1026 11
rect 912 -14 914 -6
rect 1094 -5 1096 11
rect 1102 -5 1104 11
rect 1058 -14 1060 -6
rect 2009 -5 2011 11
rect 2017 -5 2019 11
rect 1977 -14 1979 -6
rect 2087 -5 2089 11
rect 2095 -5 2097 11
rect 2155 -5 2157 11
rect 2163 -5 2165 11
rect 2051 -14 2053 -6
rect 2233 -5 2235 11
rect 2241 -5 2243 11
rect 2276 1 2278 9
rect 2197 -14 2199 -6
rect 2307 -5 2309 11
rect 2315 -5 2317 11
rect 2385 -5 2387 11
rect 2393 -5 2395 11
rect 2453 -5 2455 11
rect 2461 -5 2463 11
rect 2349 -14 2351 -6
rect 2531 -5 2533 11
rect 2539 -5 2541 11
rect 2495 -14 2497 -6
<< ndiffusion >>
rect 1970 183 1971 187
rect 1973 183 1974 187
rect 2043 168 2044 172
rect 2046 168 2047 172
rect 2189 168 2190 172
rect 2192 168 2193 172
rect 2001 154 2002 162
rect 2004 154 2005 162
rect 2009 154 2010 162
rect 2012 154 2013 162
rect 2079 154 2080 162
rect 2082 154 2083 162
rect 2087 154 2088 162
rect 2090 154 2091 162
rect 2147 154 2148 162
rect 2150 154 2151 162
rect 2155 154 2156 162
rect 2158 154 2159 162
rect 2225 154 2226 162
rect 2228 154 2229 162
rect 2233 154 2234 162
rect 2236 154 2237 162
rect -57 71 -56 75
rect -54 71 -53 75
rect 17 71 18 75
rect 20 71 21 75
rect 163 71 164 75
rect 166 71 167 75
rect 243 71 244 75
rect 246 71 247 75
rect 315 71 316 75
rect 318 71 319 75
rect 461 71 462 75
rect 464 71 465 75
rect 541 71 542 75
rect 544 71 545 75
rect 613 71 614 75
rect 616 71 617 75
rect 759 71 760 75
rect 762 71 763 75
rect 839 71 840 75
rect 842 71 843 75
rect 911 71 912 75
rect 914 71 915 75
rect 1057 71 1058 75
rect 1060 71 1061 75
rect 1976 71 1977 75
rect 1979 71 1980 75
rect 2050 71 2051 75
rect 2053 71 2054 75
rect 2196 71 2197 75
rect 2199 71 2200 75
rect 2276 71 2277 75
rect 2279 71 2280 75
rect 2348 71 2349 75
rect 2351 71 2352 75
rect 2494 71 2495 75
rect 2497 71 2498 75
rect -25 57 -24 65
rect -22 57 -21 65
rect -17 57 -16 65
rect -14 57 -13 65
rect 53 57 54 65
rect 56 57 57 65
rect 61 57 62 65
rect 64 57 65 65
rect 121 57 122 65
rect 124 57 125 65
rect 129 57 130 65
rect 132 57 133 65
rect 199 57 200 65
rect 202 57 203 65
rect 207 57 208 65
rect 210 57 211 65
rect 273 57 274 65
rect 276 57 277 65
rect 281 57 282 65
rect 284 57 285 65
rect 351 57 352 65
rect 354 57 355 65
rect 359 57 360 65
rect 362 57 363 65
rect 419 57 420 65
rect 422 57 423 65
rect 427 57 428 65
rect 430 57 431 65
rect 497 57 498 65
rect 500 57 501 65
rect 505 57 506 65
rect 508 57 509 65
rect 571 57 572 65
rect 574 57 575 65
rect 579 57 580 65
rect 582 57 583 65
rect 649 57 650 65
rect 652 57 653 65
rect 657 57 658 65
rect 660 57 661 65
rect 717 57 718 65
rect 720 57 721 65
rect 725 57 726 65
rect 728 57 729 65
rect 795 57 796 65
rect 798 57 799 65
rect 803 57 804 65
rect 806 57 807 65
rect 869 57 870 65
rect 872 57 873 65
rect 877 57 878 65
rect 880 57 881 65
rect 947 57 948 65
rect 950 57 951 65
rect 955 57 956 65
rect 958 57 959 65
rect 1015 57 1016 65
rect 1018 57 1019 65
rect 1023 57 1024 65
rect 1026 57 1027 65
rect 1093 57 1094 65
rect 1096 57 1097 65
rect 1101 57 1102 65
rect 1104 57 1105 65
rect 2008 57 2009 65
rect 2011 57 2012 65
rect 2016 57 2017 65
rect 2019 57 2020 65
rect 2086 57 2087 65
rect 2089 57 2090 65
rect 2094 57 2095 65
rect 2097 57 2098 65
rect 2154 57 2155 65
rect 2157 57 2158 65
rect 2162 57 2163 65
rect 2165 57 2166 65
rect 2232 57 2233 65
rect 2235 57 2236 65
rect 2240 57 2241 65
rect 2243 57 2244 65
rect 2306 57 2307 65
rect 2309 57 2310 65
rect 2314 57 2315 65
rect 2317 57 2318 65
rect 2384 57 2385 65
rect 2387 57 2388 65
rect 2392 57 2393 65
rect 2395 57 2396 65
rect 2452 57 2453 65
rect 2455 57 2456 65
rect 2460 57 2461 65
rect 2463 57 2464 65
rect 2530 57 2531 65
rect 2533 57 2534 65
rect 2538 57 2539 65
rect 2541 57 2542 65
rect -57 -30 -56 -26
rect -54 -30 -53 -26
rect 13 -30 18 -26
rect 20 -30 25 -26
rect 163 -30 164 -26
rect 166 -30 167 -26
rect 242 -15 243 -11
rect 245 -15 246 -11
rect 315 -30 316 -26
rect 318 -30 319 -26
rect 461 -30 462 -26
rect 464 -30 465 -26
rect 540 -15 541 -11
rect 543 -15 544 -11
rect 613 -30 614 -26
rect 616 -30 617 -26
rect 759 -30 760 -26
rect 762 -30 763 -26
rect 838 -15 839 -11
rect 841 -15 842 -11
rect 911 -30 912 -26
rect 914 -30 915 -26
rect 1057 -30 1058 -26
rect 1060 -30 1061 -26
rect 1976 -30 1977 -26
rect 1979 -30 1980 -26
rect 2050 -30 2051 -26
rect 2053 -30 2054 -26
rect 2196 -30 2197 -26
rect 2199 -30 2200 -26
rect 2275 -15 2276 -11
rect 2278 -15 2279 -11
rect 2348 -30 2349 -26
rect 2351 -30 2352 -26
rect 2494 -30 2495 -26
rect 2497 -30 2498 -26
rect -25 -44 -24 -36
rect -22 -44 -21 -36
rect -17 -44 -16 -36
rect -14 -44 -13 -36
rect 53 -44 54 -36
rect 56 -44 57 -36
rect 61 -44 62 -36
rect 64 -44 65 -36
rect 121 -44 122 -36
rect 124 -44 125 -36
rect 129 -44 130 -36
rect 132 -44 133 -36
rect 199 -44 200 -36
rect 202 -44 203 -36
rect 207 -44 208 -36
rect 210 -44 211 -36
rect 273 -44 274 -36
rect 276 -44 277 -36
rect 281 -44 282 -36
rect 284 -44 285 -36
rect 351 -44 352 -36
rect 354 -44 355 -36
rect 359 -44 360 -36
rect 362 -44 363 -36
rect 419 -44 420 -36
rect 422 -44 423 -36
rect 427 -44 428 -36
rect 430 -44 431 -36
rect 497 -44 498 -36
rect 500 -44 501 -36
rect 505 -44 506 -36
rect 508 -44 509 -36
rect 571 -44 572 -36
rect 574 -44 575 -36
rect 579 -44 580 -36
rect 582 -44 583 -36
rect 649 -44 650 -36
rect 652 -44 653 -36
rect 657 -44 658 -36
rect 660 -44 661 -36
rect 717 -44 718 -36
rect 720 -44 721 -36
rect 725 -44 726 -36
rect 728 -44 729 -36
rect 795 -44 796 -36
rect 798 -44 799 -36
rect 803 -44 804 -36
rect 806 -44 807 -36
rect 869 -44 870 -36
rect 872 -44 873 -36
rect 877 -44 878 -36
rect 880 -44 881 -36
rect 947 -44 948 -36
rect 950 -44 951 -36
rect 955 -44 956 -36
rect 958 -44 959 -36
rect 1015 -44 1016 -36
rect 1018 -44 1019 -36
rect 1023 -44 1024 -36
rect 1026 -44 1027 -36
rect 1093 -44 1094 -36
rect 1096 -44 1097 -36
rect 1101 -44 1102 -36
rect 1104 -44 1105 -36
rect 2008 -44 2009 -36
rect 2011 -44 2012 -36
rect 2016 -44 2017 -36
rect 2019 -44 2020 -36
rect 2086 -44 2087 -36
rect 2089 -44 2090 -36
rect 2094 -44 2095 -36
rect 2097 -44 2098 -36
rect 2154 -44 2155 -36
rect 2157 -44 2158 -36
rect 2162 -44 2163 -36
rect 2165 -44 2166 -36
rect 2232 -44 2233 -36
rect 2235 -44 2236 -36
rect 2240 -44 2241 -36
rect 2243 -44 2244 -36
rect 2306 -44 2307 -36
rect 2309 -44 2310 -36
rect 2314 -44 2315 -36
rect 2317 -44 2318 -36
rect 2384 -44 2385 -36
rect 2387 -44 2388 -36
rect 2392 -44 2393 -36
rect 2395 -44 2396 -36
rect 2452 -44 2453 -36
rect 2455 -44 2456 -36
rect 2460 -44 2461 -36
rect 2463 -44 2464 -36
rect 2530 -44 2531 -36
rect 2533 -44 2534 -36
rect 2538 -44 2539 -36
rect 2541 -44 2542 -36
<< pdiffusion >>
rect 1970 199 1971 207
rect 1973 199 1974 207
rect 2001 193 2002 209
rect 2004 193 2005 209
rect 2009 193 2010 209
rect 2012 193 2013 209
rect 2079 193 2080 209
rect 2082 193 2083 209
rect 2087 193 2088 209
rect 2090 193 2091 209
rect 2147 193 2148 209
rect 2150 193 2151 209
rect 2155 193 2156 209
rect 2158 193 2159 209
rect 2043 184 2044 192
rect 2046 184 2047 192
rect 2225 193 2226 209
rect 2228 193 2229 209
rect 2233 193 2234 209
rect 2236 193 2237 209
rect 2189 184 2190 192
rect 2192 184 2193 192
rect -25 96 -24 112
rect -22 96 -21 112
rect -17 96 -16 112
rect -14 96 -13 112
rect -57 87 -56 95
rect -54 87 -53 95
rect 53 96 54 112
rect 56 96 57 112
rect 61 96 62 112
rect 64 96 65 112
rect 121 96 122 112
rect 124 96 125 112
rect 129 96 130 112
rect 132 96 133 112
rect 17 87 18 95
rect 20 87 21 95
rect 199 96 200 112
rect 202 96 203 112
rect 207 96 208 112
rect 210 96 211 112
rect 163 87 164 95
rect 166 87 167 95
rect 273 96 274 112
rect 276 96 277 112
rect 281 96 282 112
rect 284 96 285 112
rect 243 87 244 95
rect 246 87 247 95
rect 351 96 352 112
rect 354 96 355 112
rect 359 96 360 112
rect 362 96 363 112
rect 419 96 420 112
rect 422 96 423 112
rect 427 96 428 112
rect 430 96 431 112
rect 315 87 316 95
rect 318 87 319 95
rect 497 96 498 112
rect 500 96 501 112
rect 505 96 506 112
rect 508 96 509 112
rect 461 87 462 95
rect 464 87 465 95
rect 571 96 572 112
rect 574 96 575 112
rect 579 96 580 112
rect 582 96 583 112
rect 541 87 542 95
rect 544 87 545 95
rect 649 96 650 112
rect 652 96 653 112
rect 657 96 658 112
rect 660 96 661 112
rect 717 96 718 112
rect 720 96 721 112
rect 725 96 726 112
rect 728 96 729 112
rect 613 87 614 95
rect 616 87 617 95
rect 795 96 796 112
rect 798 96 799 112
rect 803 96 804 112
rect 806 96 807 112
rect 759 87 760 95
rect 762 87 763 95
rect 869 96 870 112
rect 872 96 873 112
rect 877 96 878 112
rect 880 96 881 112
rect 839 87 840 95
rect 842 87 843 95
rect 947 96 948 112
rect 950 96 951 112
rect 955 96 956 112
rect 958 96 959 112
rect 1015 96 1016 112
rect 1018 96 1019 112
rect 1023 96 1024 112
rect 1026 96 1027 112
rect 911 87 912 95
rect 914 87 915 95
rect 1093 96 1094 112
rect 1096 96 1097 112
rect 1101 96 1102 112
rect 1104 96 1105 112
rect 1057 87 1058 95
rect 1060 87 1061 95
rect 2008 96 2009 112
rect 2011 96 2012 112
rect 2016 96 2017 112
rect 2019 96 2020 112
rect 1976 87 1977 95
rect 1979 87 1980 95
rect 2086 96 2087 112
rect 2089 96 2090 112
rect 2094 96 2095 112
rect 2097 96 2098 112
rect 2154 96 2155 112
rect 2157 96 2158 112
rect 2162 96 2163 112
rect 2165 96 2166 112
rect 2050 87 2051 95
rect 2053 87 2054 95
rect 2232 96 2233 112
rect 2235 96 2236 112
rect 2240 96 2241 112
rect 2243 96 2244 112
rect 2196 87 2197 95
rect 2199 87 2200 95
rect 2306 96 2307 112
rect 2309 96 2310 112
rect 2314 96 2315 112
rect 2317 96 2318 112
rect 2276 87 2277 95
rect 2279 87 2280 95
rect 2384 96 2385 112
rect 2387 96 2388 112
rect 2392 96 2393 112
rect 2395 96 2396 112
rect 2452 96 2453 112
rect 2455 96 2456 112
rect 2460 96 2461 112
rect 2463 96 2464 112
rect 2348 87 2349 95
rect 2351 87 2352 95
rect 2530 96 2531 112
rect 2533 96 2534 112
rect 2538 96 2539 112
rect 2541 96 2542 112
rect 2494 87 2495 95
rect 2497 87 2498 95
rect -25 -5 -24 11
rect -22 -5 -21 11
rect -17 -5 -16 11
rect -14 -5 -13 11
rect -57 -14 -56 -6
rect -54 -14 -53 -6
rect 53 -5 54 11
rect 56 -5 57 11
rect 61 -5 62 11
rect 64 -5 65 11
rect 121 -5 122 11
rect 124 -5 125 11
rect 129 -5 130 11
rect 132 -5 133 11
rect 13 -14 18 -6
rect 20 -14 25 -6
rect 199 -5 200 11
rect 202 -5 203 11
rect 207 -5 208 11
rect 210 -5 211 11
rect 242 1 243 9
rect 245 1 246 9
rect 163 -14 164 -6
rect 166 -14 167 -6
rect 273 -5 274 11
rect 276 -5 277 11
rect 281 -5 282 11
rect 284 -5 285 11
rect 351 -5 352 11
rect 354 -5 355 11
rect 359 -5 360 11
rect 362 -5 363 11
rect 419 -5 420 11
rect 422 -5 423 11
rect 427 -5 428 11
rect 430 -5 431 11
rect 315 -14 316 -6
rect 318 -14 319 -6
rect 497 -5 498 11
rect 500 -5 501 11
rect 505 -5 506 11
rect 508 -5 509 11
rect 540 1 541 9
rect 543 1 544 9
rect 461 -14 462 -6
rect 464 -14 465 -6
rect 571 -5 572 11
rect 574 -5 575 11
rect 579 -5 580 11
rect 582 -5 583 11
rect 649 -5 650 11
rect 652 -5 653 11
rect 657 -5 658 11
rect 660 -5 661 11
rect 717 -5 718 11
rect 720 -5 721 11
rect 725 -5 726 11
rect 728 -5 729 11
rect 613 -14 614 -6
rect 616 -14 617 -6
rect 795 -5 796 11
rect 798 -5 799 11
rect 803 -5 804 11
rect 806 -5 807 11
rect 838 1 839 9
rect 841 1 842 9
rect 759 -14 760 -6
rect 762 -14 763 -6
rect 869 -5 870 11
rect 872 -5 873 11
rect 877 -5 878 11
rect 880 -5 881 11
rect 947 -5 948 11
rect 950 -5 951 11
rect 955 -5 956 11
rect 958 -5 959 11
rect 1015 -5 1016 11
rect 1018 -5 1019 11
rect 1023 -5 1024 11
rect 1026 -5 1027 11
rect 911 -14 912 -6
rect 914 -14 915 -6
rect 1093 -5 1094 11
rect 1096 -5 1097 11
rect 1101 -5 1102 11
rect 1104 -5 1105 11
rect 1057 -14 1058 -6
rect 1060 -14 1061 -6
rect 2008 -5 2009 11
rect 2011 -5 2012 11
rect 2016 -5 2017 11
rect 2019 -5 2020 11
rect 1976 -14 1977 -6
rect 1979 -14 1980 -6
rect 2086 -5 2087 11
rect 2089 -5 2090 11
rect 2094 -5 2095 11
rect 2097 -5 2098 11
rect 2154 -5 2155 11
rect 2157 -5 2158 11
rect 2162 -5 2163 11
rect 2165 -5 2166 11
rect 2050 -14 2051 -6
rect 2053 -14 2054 -6
rect 2232 -5 2233 11
rect 2235 -5 2236 11
rect 2240 -5 2241 11
rect 2243 -5 2244 11
rect 2275 1 2276 9
rect 2278 1 2279 9
rect 2196 -14 2197 -6
rect 2199 -14 2200 -6
rect 2306 -5 2307 11
rect 2309 -5 2310 11
rect 2314 -5 2315 11
rect 2317 -5 2318 11
rect 2384 -5 2385 11
rect 2387 -5 2388 11
rect 2392 -5 2393 11
rect 2395 -5 2396 11
rect 2452 -5 2453 11
rect 2455 -5 2456 11
rect 2460 -5 2461 11
rect 2463 -5 2464 11
rect 2348 -14 2349 -6
rect 2351 -14 2352 -6
rect 2530 -5 2531 11
rect 2533 -5 2534 11
rect 2538 -5 2539 11
rect 2541 -5 2542 11
rect 2494 -14 2495 -6
rect 2497 -14 2498 -6
<< ndcontact >>
rect 1966 183 1970 187
rect 1974 183 1978 187
rect 2039 168 2043 172
rect 2047 168 2051 172
rect 2185 168 2189 172
rect 2193 168 2197 172
rect 1997 154 2001 162
rect 2005 154 2009 162
rect 2013 154 2017 162
rect 2075 154 2079 162
rect 2083 154 2087 162
rect 2091 154 2095 162
rect 2143 154 2147 162
rect 2151 154 2155 162
rect 2159 154 2163 162
rect 2221 154 2225 162
rect 2229 154 2233 162
rect 2237 154 2241 162
rect -61 71 -57 75
rect -53 71 -49 75
rect 13 71 17 75
rect 21 71 25 75
rect 159 71 163 75
rect 167 71 171 75
rect 239 71 243 75
rect 247 71 251 75
rect 311 71 315 75
rect 319 71 323 75
rect 457 71 461 75
rect 465 71 469 75
rect 537 71 541 75
rect 545 71 549 75
rect 609 71 613 75
rect 617 71 621 75
rect 755 71 759 75
rect 763 71 767 75
rect 835 71 839 75
rect 843 71 847 75
rect 907 71 911 75
rect 915 71 919 75
rect 1053 71 1057 75
rect 1061 71 1065 75
rect 1972 71 1976 75
rect 1980 71 1984 75
rect 2046 71 2050 75
rect 2054 71 2058 75
rect 2192 71 2196 75
rect 2200 71 2204 75
rect 2272 71 2276 75
rect 2280 71 2284 75
rect 2344 71 2348 75
rect 2352 71 2356 75
rect 2490 71 2494 75
rect 2498 71 2502 75
rect -29 57 -25 65
rect -21 57 -17 65
rect -13 57 -9 65
rect 49 57 53 65
rect 57 57 61 65
rect 65 57 69 65
rect 117 57 121 65
rect 125 57 129 65
rect 133 57 137 65
rect 195 57 199 65
rect 203 57 207 65
rect 211 57 215 65
rect 269 57 273 65
rect 277 57 281 65
rect 285 57 289 65
rect 347 57 351 65
rect 355 57 359 65
rect 363 57 367 65
rect 415 57 419 65
rect 423 57 427 65
rect 431 57 435 65
rect 493 57 497 65
rect 501 57 505 65
rect 509 57 513 65
rect 567 57 571 65
rect 575 57 579 65
rect 583 57 587 65
rect 645 57 649 65
rect 653 57 657 65
rect 661 57 665 65
rect 713 57 717 65
rect 721 57 725 65
rect 729 57 733 65
rect 791 57 795 65
rect 799 57 803 65
rect 807 57 811 65
rect 865 57 869 65
rect 873 57 877 65
rect 881 57 885 65
rect 943 57 947 65
rect 951 57 955 65
rect 959 57 963 65
rect 1011 57 1015 65
rect 1019 57 1023 65
rect 1027 57 1031 65
rect 1089 57 1093 65
rect 1097 57 1101 65
rect 1105 57 1109 65
rect 2004 57 2008 65
rect 2012 57 2016 65
rect 2020 57 2024 65
rect 2082 57 2086 65
rect 2090 57 2094 65
rect 2098 57 2102 65
rect 2150 57 2154 65
rect 2158 57 2162 65
rect 2166 57 2170 65
rect 2228 57 2232 65
rect 2236 57 2240 65
rect 2244 57 2248 65
rect 2302 57 2306 65
rect 2310 57 2314 65
rect 2318 57 2322 65
rect 2380 57 2384 65
rect 2388 57 2392 65
rect 2396 57 2400 65
rect 2448 57 2452 65
rect 2456 57 2460 65
rect 2464 57 2468 65
rect 2526 57 2530 65
rect 2534 57 2538 65
rect 2542 57 2546 65
rect -61 -30 -57 -26
rect -53 -30 -49 -26
rect 159 -30 163 -26
rect 167 -30 171 -26
rect 238 -15 242 -11
rect 246 -15 250 -11
rect 311 -30 315 -26
rect 319 -30 323 -26
rect 457 -30 461 -26
rect 465 -30 469 -26
rect 536 -15 540 -11
rect 544 -15 548 -11
rect 609 -30 613 -26
rect 617 -30 621 -26
rect 755 -30 759 -26
rect 763 -30 767 -26
rect 834 -15 838 -11
rect 842 -15 846 -11
rect 907 -30 911 -26
rect 915 -30 919 -26
rect 1053 -30 1057 -26
rect 1061 -30 1065 -26
rect 1972 -30 1976 -26
rect 1980 -30 1984 -26
rect 2046 -30 2050 -26
rect 2054 -30 2058 -26
rect 2192 -30 2196 -26
rect 2200 -30 2204 -26
rect 2271 -15 2275 -11
rect 2279 -15 2283 -11
rect 2344 -30 2348 -26
rect 2352 -30 2356 -26
rect 2490 -30 2494 -26
rect 2498 -30 2502 -26
rect -29 -44 -25 -36
rect -21 -44 -17 -36
rect -13 -44 -9 -36
rect 49 -44 53 -36
rect 57 -44 61 -36
rect 65 -44 69 -36
rect 117 -44 121 -36
rect 125 -44 129 -36
rect 133 -44 137 -36
rect 195 -44 199 -36
rect 203 -44 207 -36
rect 211 -44 215 -36
rect 269 -44 273 -36
rect 277 -44 281 -36
rect 285 -44 289 -36
rect 347 -44 351 -36
rect 355 -44 359 -36
rect 363 -44 367 -36
rect 415 -44 419 -36
rect 423 -44 427 -36
rect 431 -44 435 -36
rect 493 -44 497 -36
rect 501 -44 505 -36
rect 509 -44 513 -36
rect 567 -44 571 -36
rect 575 -44 579 -36
rect 583 -44 587 -36
rect 645 -44 649 -36
rect 653 -44 657 -36
rect 661 -44 665 -36
rect 713 -44 717 -36
rect 721 -44 725 -36
rect 729 -44 733 -36
rect 791 -44 795 -36
rect 799 -44 803 -36
rect 807 -44 811 -36
rect 865 -44 869 -36
rect 873 -44 877 -36
rect 881 -44 885 -36
rect 943 -44 947 -36
rect 951 -44 955 -36
rect 959 -44 963 -36
rect 1011 -44 1015 -36
rect 1019 -44 1023 -36
rect 1027 -44 1031 -36
rect 1089 -44 1093 -36
rect 1097 -44 1101 -36
rect 1105 -44 1109 -36
rect 2004 -44 2008 -36
rect 2012 -44 2016 -36
rect 2020 -44 2024 -36
rect 2082 -44 2086 -36
rect 2090 -44 2094 -36
rect 2098 -44 2102 -36
rect 2150 -44 2154 -36
rect 2158 -44 2162 -36
rect 2166 -44 2170 -36
rect 2228 -44 2232 -36
rect 2236 -44 2240 -36
rect 2244 -44 2248 -36
rect 2302 -44 2306 -36
rect 2310 -44 2314 -36
rect 2318 -44 2322 -36
rect 2380 -44 2384 -36
rect 2388 -44 2392 -36
rect 2396 -44 2400 -36
rect 2448 -44 2452 -36
rect 2456 -44 2460 -36
rect 2464 -44 2468 -36
rect 2526 -44 2530 -36
rect 2534 -44 2538 -36
rect 2542 -44 2546 -36
<< pdcontact >>
rect 1966 199 1970 207
rect 1974 199 1978 207
rect 1997 193 2001 209
rect 2005 193 2009 209
rect 2013 193 2017 209
rect 2075 193 2079 209
rect 2083 193 2087 209
rect 2091 193 2095 209
rect 2143 193 2147 209
rect 2151 193 2155 209
rect 2159 193 2163 209
rect 2039 184 2043 192
rect 2047 184 2051 192
rect 2221 193 2225 209
rect 2229 193 2233 209
rect 2237 193 2241 209
rect 2185 184 2189 192
rect 2193 184 2197 192
rect -29 96 -25 112
rect -21 96 -17 112
rect -13 96 -9 112
rect -61 87 -57 95
rect -53 87 -49 95
rect 49 96 53 112
rect 57 96 61 112
rect 65 96 69 112
rect 117 96 121 112
rect 125 96 129 112
rect 133 96 137 112
rect 13 87 17 95
rect 21 87 25 95
rect 195 96 199 112
rect 203 96 207 112
rect 211 96 215 112
rect 159 87 163 95
rect 167 87 171 95
rect 269 96 273 112
rect 277 96 281 112
rect 285 96 289 112
rect 239 87 243 95
rect 247 87 251 95
rect 347 96 351 112
rect 355 96 359 112
rect 363 96 367 112
rect 415 96 419 112
rect 423 96 427 112
rect 431 96 435 112
rect 311 87 315 95
rect 319 87 323 95
rect 493 96 497 112
rect 501 96 505 112
rect 509 96 513 112
rect 457 87 461 95
rect 465 87 469 95
rect 567 96 571 112
rect 575 96 579 112
rect 583 96 587 112
rect 537 87 541 95
rect 545 87 549 95
rect 645 96 649 112
rect 653 96 657 112
rect 661 96 665 112
rect 713 96 717 112
rect 721 96 725 112
rect 729 96 733 112
rect 609 87 613 95
rect 617 87 621 95
rect 791 96 795 112
rect 799 96 803 112
rect 807 96 811 112
rect 755 87 759 95
rect 763 87 767 95
rect 865 96 869 112
rect 873 96 877 112
rect 881 96 885 112
rect 835 87 839 95
rect 843 87 847 95
rect 943 96 947 112
rect 951 96 955 112
rect 959 96 963 112
rect 1011 96 1015 112
rect 1019 96 1023 112
rect 1027 96 1031 112
rect 907 87 911 95
rect 915 87 919 95
rect 1089 96 1093 112
rect 1097 96 1101 112
rect 1105 96 1109 112
rect 1053 87 1057 95
rect 1061 87 1065 95
rect 2004 96 2008 112
rect 2012 96 2016 112
rect 2020 96 2024 112
rect 1972 87 1976 95
rect 1980 87 1984 95
rect 2082 96 2086 112
rect 2090 96 2094 112
rect 2098 96 2102 112
rect 2150 96 2154 112
rect 2158 96 2162 112
rect 2166 96 2170 112
rect 2046 87 2050 95
rect 2054 87 2058 95
rect 2228 96 2232 112
rect 2236 96 2240 112
rect 2244 96 2248 112
rect 2192 87 2196 95
rect 2200 87 2204 95
rect 2302 96 2306 112
rect 2310 96 2314 112
rect 2318 96 2322 112
rect 2272 87 2276 95
rect 2280 87 2284 95
rect 2380 96 2384 112
rect 2388 96 2392 112
rect 2396 96 2400 112
rect 2448 96 2452 112
rect 2456 96 2460 112
rect 2464 96 2468 112
rect 2344 87 2348 95
rect 2352 87 2356 95
rect 2526 96 2530 112
rect 2534 96 2538 112
rect 2542 96 2546 112
rect 2490 87 2494 95
rect 2498 87 2502 95
rect -29 -5 -25 11
rect -21 -5 -17 11
rect -13 -5 -9 11
rect -61 -14 -57 -6
rect -53 -14 -49 -6
rect 49 -5 53 11
rect 57 -5 61 11
rect 65 -5 69 11
rect 117 -5 121 11
rect 125 -5 129 11
rect 133 -5 137 11
rect 195 -5 199 11
rect 203 -5 207 11
rect 211 -5 215 11
rect 238 1 242 9
rect 246 1 250 9
rect 159 -14 163 -6
rect 167 -14 171 -6
rect 269 -5 273 11
rect 277 -5 281 11
rect 285 -5 289 11
rect 347 -5 351 11
rect 355 -5 359 11
rect 363 -5 367 11
rect 415 -5 419 11
rect 423 -5 427 11
rect 431 -5 435 11
rect 311 -14 315 -6
rect 319 -14 323 -6
rect 493 -5 497 11
rect 501 -5 505 11
rect 509 -5 513 11
rect 536 1 540 9
rect 544 1 548 9
rect 457 -14 461 -6
rect 465 -14 469 -6
rect 567 -5 571 11
rect 575 -5 579 11
rect 583 -5 587 11
rect 645 -5 649 11
rect 653 -5 657 11
rect 661 -5 665 11
rect 713 -5 717 11
rect 721 -5 725 11
rect 729 -5 733 11
rect 609 -14 613 -6
rect 617 -14 621 -6
rect 791 -5 795 11
rect 799 -5 803 11
rect 807 -5 811 11
rect 834 1 838 9
rect 842 1 846 9
rect 755 -14 759 -6
rect 763 -14 767 -6
rect 865 -5 869 11
rect 873 -5 877 11
rect 881 -5 885 11
rect 943 -5 947 11
rect 951 -5 955 11
rect 959 -5 963 11
rect 1011 -5 1015 11
rect 1019 -5 1023 11
rect 1027 -5 1031 11
rect 907 -14 911 -6
rect 915 -14 919 -6
rect 1089 -5 1093 11
rect 1097 -5 1101 11
rect 1105 -5 1109 11
rect 1053 -14 1057 -6
rect 1061 -14 1065 -6
rect 2004 -5 2008 11
rect 2012 -5 2016 11
rect 2020 -5 2024 11
rect 1972 -14 1976 -6
rect 1980 -14 1984 -6
rect 2082 -5 2086 11
rect 2090 -5 2094 11
rect 2098 -5 2102 11
rect 2150 -5 2154 11
rect 2158 -5 2162 11
rect 2166 -5 2170 11
rect 2046 -14 2050 -6
rect 2054 -14 2058 -6
rect 2228 -5 2232 11
rect 2236 -5 2240 11
rect 2244 -5 2248 11
rect 2271 1 2275 9
rect 2279 1 2283 9
rect 2192 -14 2196 -6
rect 2200 -14 2204 -6
rect 2302 -5 2306 11
rect 2310 -5 2314 11
rect 2318 -5 2322 11
rect 2380 -5 2384 11
rect 2388 -5 2392 11
rect 2396 -5 2400 11
rect 2448 -5 2452 11
rect 2456 -5 2460 11
rect 2464 -5 2468 11
rect 2344 -14 2348 -6
rect 2352 -14 2356 -6
rect 2526 -5 2530 11
rect 2534 -5 2538 11
rect 2542 -5 2546 11
rect 2490 -14 2494 -6
rect 2498 -14 2502 -6
<< polysilicon >>
rect 1971 207 1973 210
rect 2002 209 2004 212
rect 2010 209 2012 212
rect 2080 209 2082 212
rect 2088 209 2090 212
rect 2148 209 2150 212
rect 2156 209 2158 212
rect 2226 209 2228 212
rect 2234 209 2236 212
rect 1971 187 1973 199
rect 1971 180 1973 183
rect 2002 162 2004 193
rect 2010 179 2012 193
rect 2044 192 2046 195
rect 2010 162 2012 176
rect 2044 172 2046 184
rect 2044 165 2046 168
rect 2080 162 2082 193
rect 2088 181 2090 193
rect 2088 162 2090 174
rect 2148 162 2150 193
rect 2156 179 2158 193
rect 2190 192 2192 195
rect 2156 162 2158 176
rect 2190 172 2192 184
rect 2190 165 2192 168
rect 2226 162 2228 193
rect 2234 181 2236 193
rect 2234 162 2236 174
rect 2002 151 2004 154
rect 2010 151 2012 154
rect 2080 151 2082 154
rect 2088 151 2090 154
rect 2148 151 2150 154
rect 2156 151 2158 154
rect 2226 151 2228 154
rect 2234 151 2236 154
rect -24 112 -22 115
rect -16 112 -14 115
rect 54 112 56 115
rect 62 112 64 115
rect 122 112 124 115
rect 130 112 132 115
rect 200 112 202 115
rect 208 112 210 115
rect 274 112 276 115
rect 282 112 284 115
rect 352 112 354 115
rect 360 112 362 115
rect 420 112 422 115
rect 428 112 430 115
rect 498 112 500 115
rect 506 112 508 115
rect 572 112 574 115
rect 580 112 582 115
rect 650 112 652 115
rect 658 112 660 115
rect 718 112 720 115
rect 726 112 728 115
rect 796 112 798 115
rect 804 112 806 115
rect 870 112 872 115
rect 878 112 880 115
rect 948 112 950 115
rect 956 112 958 115
rect 1016 112 1018 115
rect 1024 112 1026 115
rect 1094 112 1096 115
rect 1102 112 1104 115
rect 2009 112 2011 115
rect 2017 112 2019 115
rect 2087 112 2089 115
rect 2095 112 2097 115
rect 2155 112 2157 115
rect 2163 112 2165 115
rect 2233 112 2235 115
rect 2241 112 2243 115
rect 2307 112 2309 115
rect 2315 112 2317 115
rect 2385 112 2387 115
rect 2393 112 2395 115
rect 2453 112 2455 115
rect 2461 112 2463 115
rect 2531 112 2533 115
rect 2539 112 2541 115
rect -56 95 -54 98
rect -56 75 -54 87
rect -56 68 -54 71
rect -24 65 -22 96
rect -16 82 -14 96
rect 18 95 20 98
rect -16 65 -14 79
rect 18 75 20 87
rect 18 68 20 71
rect 54 65 56 96
rect 62 84 64 96
rect 62 65 64 77
rect 122 65 124 96
rect 130 82 132 96
rect 164 95 166 98
rect 130 65 132 79
rect 164 75 166 87
rect 164 68 166 71
rect 200 65 202 96
rect 208 84 210 96
rect 244 95 246 98
rect 208 65 210 77
rect 244 75 246 87
rect 244 68 246 71
rect 274 65 276 96
rect 282 82 284 96
rect 316 95 318 98
rect 282 65 284 79
rect 316 75 318 87
rect 316 68 318 71
rect 352 65 354 96
rect 360 84 362 96
rect 360 65 362 77
rect 420 65 422 96
rect 428 82 430 96
rect 462 95 464 98
rect 428 65 430 79
rect 462 75 464 87
rect 462 68 464 71
rect 498 65 500 96
rect 506 84 508 96
rect 542 95 544 98
rect 506 65 508 77
rect 542 75 544 87
rect 542 68 544 71
rect 572 65 574 96
rect 580 82 582 96
rect 614 95 616 98
rect 580 65 582 79
rect 614 75 616 87
rect 614 68 616 71
rect 650 65 652 96
rect 658 84 660 96
rect 658 65 660 77
rect 718 65 720 96
rect 726 82 728 96
rect 760 95 762 98
rect 726 65 728 79
rect 760 75 762 87
rect 760 68 762 71
rect 796 65 798 96
rect 804 84 806 96
rect 840 95 842 98
rect 804 65 806 77
rect 840 75 842 87
rect 840 68 842 71
rect 870 65 872 96
rect 878 82 880 96
rect 912 95 914 98
rect 878 65 880 79
rect 912 75 914 87
rect 912 68 914 71
rect 948 65 950 96
rect 956 84 958 96
rect 956 65 958 77
rect 1016 65 1018 96
rect 1024 82 1026 96
rect 1058 95 1060 98
rect 1024 65 1026 79
rect 1058 75 1060 87
rect 1058 68 1060 71
rect 1094 65 1096 96
rect 1102 84 1104 96
rect 1977 95 1979 98
rect 1102 65 1104 77
rect 1977 75 1979 87
rect 1977 68 1979 71
rect 2009 65 2011 96
rect 2017 82 2019 96
rect 2051 95 2053 98
rect 2017 65 2019 79
rect 2051 75 2053 87
rect 2051 68 2053 71
rect 2087 65 2089 96
rect 2095 84 2097 96
rect 2095 65 2097 77
rect 2155 65 2157 96
rect 2163 82 2165 96
rect 2197 95 2199 98
rect 2163 65 2165 79
rect 2197 75 2199 87
rect 2197 68 2199 71
rect 2233 65 2235 96
rect 2241 84 2243 96
rect 2277 95 2279 98
rect 2241 65 2243 77
rect 2277 75 2279 87
rect 2277 68 2279 71
rect 2307 65 2309 96
rect 2315 82 2317 96
rect 2349 95 2351 98
rect 2315 65 2317 79
rect 2349 75 2351 87
rect 2349 68 2351 71
rect 2385 65 2387 96
rect 2393 84 2395 96
rect 2393 65 2395 77
rect 2453 65 2455 96
rect 2461 82 2463 96
rect 2495 95 2497 98
rect 2461 65 2463 79
rect 2495 75 2497 87
rect 2495 68 2497 71
rect 2531 65 2533 96
rect 2539 84 2541 96
rect 2539 65 2541 77
rect -24 54 -22 57
rect -16 54 -14 57
rect 54 54 56 57
rect 62 54 64 57
rect 122 54 124 57
rect 130 54 132 57
rect 200 54 202 57
rect 208 54 210 57
rect 274 54 276 57
rect 282 54 284 57
rect 352 54 354 57
rect 360 54 362 57
rect 420 54 422 57
rect 428 54 430 57
rect 498 54 500 57
rect 506 54 508 57
rect 572 54 574 57
rect 580 54 582 57
rect 650 54 652 57
rect 658 54 660 57
rect 718 54 720 57
rect 726 54 728 57
rect 796 54 798 57
rect 804 54 806 57
rect 870 54 872 57
rect 878 54 880 57
rect 948 54 950 57
rect 956 54 958 57
rect 1016 54 1018 57
rect 1024 54 1026 57
rect 1094 54 1096 57
rect 1102 54 1104 57
rect 2009 54 2011 57
rect 2017 54 2019 57
rect 2087 54 2089 57
rect 2095 54 2097 57
rect 2155 54 2157 57
rect 2163 54 2165 57
rect 2233 54 2235 57
rect 2241 54 2243 57
rect 2307 54 2309 57
rect 2315 54 2317 57
rect 2385 54 2387 57
rect 2393 54 2395 57
rect 2453 54 2455 57
rect 2461 54 2463 57
rect 2531 54 2533 57
rect 2539 54 2541 57
rect -24 11 -22 14
rect -16 11 -14 14
rect 54 11 56 14
rect 62 11 64 14
rect 122 11 124 14
rect 130 11 132 14
rect 200 11 202 14
rect 208 11 210 14
rect -56 -6 -54 -3
rect -56 -26 -54 -14
rect -56 -33 -54 -30
rect -24 -36 -22 -5
rect -16 -19 -14 -5
rect 18 -6 20 -3
rect -16 -36 -14 -22
rect 18 -26 20 -14
rect 18 -33 20 -30
rect 54 -36 56 -5
rect 62 -17 64 -5
rect 62 -36 64 -24
rect 122 -36 124 -5
rect 130 -19 132 -5
rect 164 -6 166 -3
rect 243 9 245 12
rect 274 11 276 14
rect 282 11 284 14
rect 352 11 354 14
rect 360 11 362 14
rect 420 11 422 14
rect 428 11 430 14
rect 498 11 500 14
rect 506 11 508 14
rect 130 -36 132 -22
rect 164 -26 166 -14
rect 164 -33 166 -30
rect 200 -36 202 -5
rect 208 -17 210 -5
rect 243 -11 245 1
rect 243 -18 245 -15
rect 208 -36 210 -24
rect 274 -36 276 -5
rect 282 -19 284 -5
rect 316 -6 318 -3
rect 282 -36 284 -22
rect 316 -26 318 -14
rect 316 -33 318 -30
rect 352 -36 354 -5
rect 360 -17 362 -5
rect 360 -36 362 -24
rect 420 -36 422 -5
rect 428 -19 430 -5
rect 462 -6 464 -3
rect 541 9 543 12
rect 572 11 574 14
rect 580 11 582 14
rect 650 11 652 14
rect 658 11 660 14
rect 718 11 720 14
rect 726 11 728 14
rect 796 11 798 14
rect 804 11 806 14
rect 428 -36 430 -22
rect 462 -26 464 -14
rect 462 -33 464 -30
rect 498 -36 500 -5
rect 506 -17 508 -5
rect 541 -11 543 1
rect 541 -18 543 -15
rect 506 -36 508 -24
rect 572 -36 574 -5
rect 580 -19 582 -5
rect 614 -6 616 -3
rect 580 -36 582 -22
rect 614 -26 616 -14
rect 614 -33 616 -30
rect 650 -36 652 -5
rect 658 -17 660 -5
rect 658 -36 660 -24
rect 718 -36 720 -5
rect 726 -19 728 -5
rect 760 -6 762 -3
rect 839 9 841 12
rect 870 11 872 14
rect 878 11 880 14
rect 948 11 950 14
rect 956 11 958 14
rect 1016 11 1018 14
rect 1024 11 1026 14
rect 1094 11 1096 14
rect 1102 11 1104 14
rect 2009 11 2011 14
rect 2017 11 2019 14
rect 2087 11 2089 14
rect 2095 11 2097 14
rect 2155 11 2157 14
rect 2163 11 2165 14
rect 2233 11 2235 14
rect 2241 11 2243 14
rect 726 -36 728 -22
rect 760 -26 762 -14
rect 760 -33 762 -30
rect 796 -36 798 -5
rect 804 -17 806 -5
rect 839 -11 841 1
rect 839 -18 841 -15
rect 804 -36 806 -24
rect 870 -36 872 -5
rect 878 -19 880 -5
rect 912 -6 914 -3
rect 878 -36 880 -22
rect 912 -26 914 -14
rect 912 -33 914 -30
rect 948 -36 950 -5
rect 956 -17 958 -5
rect 956 -36 958 -24
rect 1016 -36 1018 -5
rect 1024 -19 1026 -5
rect 1058 -6 1060 -3
rect 1024 -36 1026 -22
rect 1058 -26 1060 -14
rect 1058 -33 1060 -30
rect 1094 -36 1096 -5
rect 1102 -17 1104 -5
rect 1977 -6 1979 -3
rect 1102 -36 1104 -24
rect 1977 -26 1979 -14
rect 1977 -33 1979 -30
rect 2009 -36 2011 -5
rect 2017 -19 2019 -5
rect 2051 -6 2053 -3
rect 2017 -36 2019 -22
rect 2051 -26 2053 -14
rect 2051 -33 2053 -30
rect 2087 -36 2089 -5
rect 2095 -17 2097 -5
rect 2095 -36 2097 -24
rect 2155 -36 2157 -5
rect 2163 -19 2165 -5
rect 2197 -6 2199 -3
rect 2276 9 2278 12
rect 2307 11 2309 14
rect 2315 11 2317 14
rect 2385 11 2387 14
rect 2393 11 2395 14
rect 2453 11 2455 14
rect 2461 11 2463 14
rect 2531 11 2533 14
rect 2539 11 2541 14
rect 2163 -36 2165 -22
rect 2197 -26 2199 -14
rect 2197 -33 2199 -30
rect 2233 -36 2235 -5
rect 2241 -17 2243 -5
rect 2276 -11 2278 1
rect 2276 -18 2278 -15
rect 2241 -36 2243 -24
rect 2307 -36 2309 -5
rect 2315 -19 2317 -5
rect 2349 -6 2351 -3
rect 2315 -36 2317 -22
rect 2349 -26 2351 -14
rect 2349 -33 2351 -30
rect 2385 -36 2387 -5
rect 2393 -17 2395 -5
rect 2393 -36 2395 -24
rect 2453 -36 2455 -5
rect 2461 -19 2463 -5
rect 2495 -6 2497 -3
rect 2461 -36 2463 -22
rect 2495 -26 2497 -14
rect 2495 -33 2497 -30
rect 2531 -36 2533 -5
rect 2539 -17 2541 -5
rect 2539 -36 2541 -24
rect -24 -47 -22 -44
rect -16 -47 -14 -44
rect 54 -47 56 -44
rect 62 -47 64 -44
rect 122 -47 124 -44
rect 130 -47 132 -44
rect 200 -47 202 -44
rect 208 -47 210 -44
rect 274 -47 276 -44
rect 282 -47 284 -44
rect 352 -47 354 -44
rect 360 -47 362 -44
rect 420 -47 422 -44
rect 428 -47 430 -44
rect 498 -47 500 -44
rect 506 -47 508 -44
rect 572 -47 574 -44
rect 580 -47 582 -44
rect 650 -47 652 -44
rect 658 -47 660 -44
rect 718 -47 720 -44
rect 726 -47 728 -44
rect 796 -47 798 -44
rect 804 -47 806 -44
rect 870 -47 872 -44
rect 878 -47 880 -44
rect 948 -47 950 -44
rect 956 -47 958 -44
rect 1016 -47 1018 -44
rect 1024 -47 1026 -44
rect 1094 -47 1096 -44
rect 1102 -47 1104 -44
rect 2009 -47 2011 -44
rect 2017 -47 2019 -44
rect 2087 -47 2089 -44
rect 2095 -47 2097 -44
rect 2155 -47 2157 -44
rect 2163 -47 2165 -44
rect 2233 -47 2235 -44
rect 2241 -47 2243 -44
rect 2307 -47 2309 -44
rect 2315 -47 2317 -44
rect 2385 -47 2387 -44
rect 2393 -47 2395 -44
rect 2453 -47 2455 -44
rect 2461 -47 2463 -44
rect 2531 -47 2533 -44
rect 2539 -47 2541 -44
<< polycontact >>
rect 1967 190 1971 194
rect 1998 175 2002 179
rect 2012 182 2016 186
rect 2040 175 2044 179
rect 2076 175 2080 179
rect 2012 168 2016 172
rect 2090 182 2094 186
rect 2144 175 2148 179
rect 2090 168 2094 172
rect 2158 182 2162 186
rect 2186 175 2190 179
rect 2222 175 2226 179
rect 2158 168 2162 172
rect 2236 182 2240 186
rect 2236 168 2240 172
rect -60 78 -56 82
rect -28 78 -24 82
rect -14 85 -10 89
rect 14 78 18 82
rect 50 78 54 82
rect -14 71 -10 75
rect 64 85 68 89
rect 118 78 122 82
rect 64 71 68 75
rect 132 85 136 89
rect 160 78 164 82
rect 196 78 200 82
rect 132 71 136 75
rect 210 85 214 89
rect 240 78 244 82
rect 270 78 274 82
rect 210 71 214 75
rect 284 85 288 89
rect 312 78 316 82
rect 348 78 352 82
rect 284 71 288 75
rect 362 85 366 89
rect 416 78 420 82
rect 362 71 366 75
rect 430 85 434 89
rect 458 78 462 82
rect 494 78 498 82
rect 430 71 434 75
rect 508 85 512 89
rect 538 78 542 82
rect 568 78 572 82
rect 508 71 512 75
rect 582 85 586 89
rect 610 78 614 82
rect 646 78 650 82
rect 582 71 586 75
rect 660 85 664 89
rect 714 78 718 82
rect 660 71 664 75
rect 728 85 732 89
rect 756 78 760 82
rect 792 78 796 82
rect 728 71 732 75
rect 806 85 810 89
rect 836 78 840 82
rect 866 78 870 82
rect 806 71 810 75
rect 880 85 884 89
rect 908 78 912 82
rect 944 78 948 82
rect 880 71 884 75
rect 958 85 962 89
rect 1012 78 1016 82
rect 958 71 962 75
rect 1026 85 1030 89
rect 1054 78 1058 82
rect 1090 78 1094 82
rect 1026 71 1030 75
rect 1104 85 1108 89
rect 1973 78 1977 82
rect 2005 78 2009 82
rect 1104 71 1108 75
rect 2019 85 2023 89
rect 2047 78 2051 82
rect 2083 78 2087 82
rect 2019 71 2023 75
rect 2097 85 2101 89
rect 2151 78 2155 82
rect 2097 71 2101 75
rect 2165 85 2169 89
rect 2193 78 2197 82
rect 2229 78 2233 82
rect 2165 71 2169 75
rect 2243 85 2247 89
rect 2273 78 2277 82
rect 2303 78 2307 82
rect 2243 71 2247 75
rect 2317 85 2321 89
rect 2345 78 2349 82
rect 2381 78 2385 82
rect 2317 71 2321 75
rect 2395 85 2399 89
rect 2449 78 2453 82
rect 2395 71 2399 75
rect 2463 85 2467 89
rect 2491 78 2495 82
rect 2527 78 2531 82
rect 2463 71 2467 75
rect 2541 85 2545 89
rect 2541 71 2545 75
rect -60 -23 -56 -19
rect -28 -23 -24 -19
rect -14 -16 -10 -12
rect 14 -23 18 -19
rect 50 -23 54 -19
rect -14 -30 -10 -26
rect 64 -16 68 -12
rect 118 -23 122 -19
rect 64 -30 68 -26
rect 132 -16 136 -12
rect 160 -23 164 -19
rect 196 -23 200 -19
rect 132 -30 136 -26
rect 239 -8 243 -4
rect 210 -16 214 -12
rect 270 -23 274 -19
rect 210 -30 214 -26
rect 284 -16 288 -12
rect 312 -23 316 -19
rect 348 -23 352 -19
rect 284 -30 288 -26
rect 362 -16 366 -12
rect 416 -23 420 -19
rect 362 -30 366 -26
rect 430 -16 434 -12
rect 458 -23 462 -19
rect 494 -23 498 -19
rect 430 -30 434 -26
rect 537 -8 541 -4
rect 508 -16 512 -12
rect 568 -23 572 -19
rect 508 -30 512 -26
rect 582 -16 586 -12
rect 610 -23 614 -19
rect 646 -23 650 -19
rect 582 -30 586 -26
rect 660 -16 664 -12
rect 714 -23 718 -19
rect 660 -30 664 -26
rect 728 -16 732 -12
rect 756 -23 760 -19
rect 792 -23 796 -19
rect 728 -30 732 -26
rect 835 -8 839 -4
rect 806 -16 810 -12
rect 866 -23 870 -19
rect 806 -30 810 -26
rect 880 -16 884 -12
rect 908 -23 912 -19
rect 944 -23 948 -19
rect 880 -30 884 -26
rect 958 -16 962 -12
rect 1012 -23 1016 -19
rect 958 -30 962 -26
rect 1026 -16 1030 -12
rect 1054 -23 1058 -19
rect 1090 -23 1094 -19
rect 1026 -30 1030 -26
rect 1104 -16 1108 -12
rect 1973 -23 1977 -19
rect 2005 -23 2009 -19
rect 1104 -30 1108 -26
rect 2019 -16 2023 -12
rect 2047 -23 2051 -19
rect 2083 -23 2087 -19
rect 2019 -30 2023 -26
rect 2097 -16 2101 -12
rect 2151 -23 2155 -19
rect 2097 -30 2101 -26
rect 2165 -16 2169 -12
rect 2193 -23 2197 -19
rect 2229 -23 2233 -19
rect 2165 -30 2169 -26
rect 2272 -8 2276 -4
rect 2243 -16 2247 -12
rect 2303 -23 2307 -19
rect 2243 -30 2247 -26
rect 2317 -16 2321 -12
rect 2345 -23 2349 -19
rect 2381 -23 2385 -19
rect 2317 -30 2321 -26
rect 2395 -16 2399 -12
rect 2449 -23 2453 -19
rect 2395 -30 2399 -26
rect 2463 -16 2467 -12
rect 2491 -23 2495 -19
rect 2527 -23 2531 -19
rect 2463 -30 2467 -26
rect 2541 -16 2545 -12
rect 2541 -30 2545 -26
<< metal1 >>
rect 1966 213 2285 216
rect 1966 207 1970 213
rect 1997 209 2001 213
rect 1964 190 1967 194
rect 1974 187 1978 199
rect 2039 199 2043 213
rect 2075 209 2079 213
rect 2143 209 2147 213
rect 2033 196 2057 199
rect 234 161 1131 165
rect 532 153 1131 157
rect 1966 150 1970 183
rect 2013 190 2023 193
rect 1974 172 1978 183
rect 1986 182 2012 186
rect 2020 179 2023 190
rect 2039 192 2043 196
rect 2047 179 2051 184
rect 2060 179 2064 206
rect 2185 199 2189 213
rect 2221 209 2225 213
rect 2179 196 2203 199
rect 2091 190 2100 193
rect 2074 182 2090 186
rect 1986 175 1998 179
rect 2020 175 2040 179
rect 2047 175 2076 179
rect 1974 168 2012 172
rect 2020 165 2023 175
rect 2047 172 2051 175
rect 2013 162 2023 165
rect 2039 164 2043 168
rect 2077 168 2090 172
rect 2097 165 2100 190
rect 2159 190 2169 193
rect 2131 182 2158 186
rect 2166 179 2169 190
rect 2185 192 2189 196
rect 2193 179 2197 184
rect 2206 179 2210 206
rect 2237 190 2246 193
rect 2220 182 2236 186
rect 2108 175 2144 179
rect 2166 175 2186 179
rect 2193 175 2222 179
rect 2127 168 2158 172
rect 2033 161 2057 164
rect 2091 162 2100 165
rect 2166 165 2169 175
rect 2193 172 2197 175
rect 2159 162 2169 165
rect 2185 164 2189 168
rect 2223 168 2236 172
rect 2243 165 2246 190
rect 2260 171 2272 175
rect 1997 150 2001 154
rect 2039 150 2043 161
rect 2179 161 2203 164
rect 2237 162 2246 165
rect 2075 150 2079 154
rect 2143 150 2147 154
rect 2185 150 2189 161
rect 2281 156 2285 213
rect 2221 150 2225 154
rect 830 145 1131 149
rect 1948 147 2225 150
rect 2254 152 2285 156
rect 1128 137 1131 141
rect 1948 119 1952 147
rect 2254 119 2258 152
rect 2267 137 2576 141
rect 2521 123 2577 127
rect -77 116 2577 119
rect -85 -48 -81 50
rect -77 18 -73 116
rect -61 95 -57 116
rect -29 112 -25 116
rect 13 102 17 116
rect 49 112 53 116
rect 117 112 121 116
rect 7 99 31 102
rect -13 93 -3 96
rect -64 78 -60 82
rect -53 75 -49 87
rect -40 85 -14 89
rect -6 82 -3 93
rect 13 95 17 99
rect 21 82 25 87
rect 34 82 38 109
rect 159 102 163 116
rect 195 112 199 116
rect 153 99 177 102
rect 65 93 74 96
rect 48 85 64 89
rect -40 78 -28 82
rect -6 78 14 82
rect 21 78 50 82
rect -49 71 -14 75
rect -61 54 -57 71
rect -6 68 -3 78
rect 21 75 25 78
rect -13 65 -3 68
rect 13 67 17 71
rect 51 71 64 75
rect 71 68 74 93
rect 133 93 143 96
rect 105 85 132 89
rect 140 82 143 93
rect 159 95 163 99
rect 167 82 171 87
rect 180 82 184 109
rect 211 93 220 96
rect 194 85 210 89
rect 82 78 118 82
rect 140 78 160 82
rect 167 78 196 82
rect 101 71 132 75
rect -65 53 -57 54
rect 7 64 31 67
rect 65 65 74 68
rect 140 68 143 78
rect 167 75 171 78
rect 133 65 143 68
rect 159 67 163 71
rect 197 71 210 75
rect 217 68 220 93
rect 239 95 243 116
rect 269 112 273 116
rect 311 102 315 116
rect 347 112 351 116
rect 415 112 419 116
rect 305 99 329 102
rect 285 93 295 96
rect 237 78 240 82
rect 247 75 251 87
rect 258 85 284 89
rect 292 82 295 93
rect 311 95 315 99
rect 319 82 323 87
rect 332 82 336 109
rect 457 102 461 116
rect 493 112 497 116
rect 451 99 475 102
rect 363 93 372 96
rect 346 85 362 89
rect 258 78 270 82
rect 292 78 312 82
rect 319 78 348 82
rect 251 71 284 75
rect -29 53 -25 57
rect 13 53 17 64
rect 153 64 177 67
rect 211 65 220 68
rect 49 53 53 57
rect 117 53 121 57
rect 159 53 163 64
rect 195 53 199 57
rect 239 53 243 71
rect 292 68 295 78
rect 319 75 323 78
rect 285 65 295 68
rect 311 67 315 71
rect 349 71 362 75
rect 369 68 372 93
rect 431 93 441 96
rect 403 85 430 89
rect 438 82 441 93
rect 457 95 461 99
rect 465 82 469 87
rect 478 82 482 109
rect 509 93 518 96
rect 492 85 508 89
rect 380 78 416 82
rect 438 78 458 82
rect 465 78 494 82
rect 399 71 430 75
rect 305 64 329 67
rect 363 65 372 68
rect 438 68 441 78
rect 465 75 469 78
rect 431 65 441 68
rect 457 67 461 71
rect 495 71 508 75
rect 515 68 518 93
rect 537 95 541 116
rect 567 112 571 116
rect 609 102 613 116
rect 645 112 649 116
rect 713 112 717 116
rect 603 99 627 102
rect 583 93 593 96
rect 535 78 538 82
rect 545 75 549 87
rect 556 85 582 89
rect 590 82 593 93
rect 609 95 613 99
rect 617 82 621 87
rect 630 82 634 109
rect 755 102 759 116
rect 791 112 795 116
rect 749 99 773 102
rect 661 93 670 96
rect 644 85 660 89
rect 556 78 568 82
rect 590 78 610 82
rect 617 78 646 82
rect 549 71 582 75
rect 269 53 273 57
rect 311 53 315 64
rect 451 64 475 67
rect 509 65 518 68
rect 347 53 351 57
rect 415 53 419 57
rect 457 53 461 64
rect 493 53 497 57
rect 537 53 541 71
rect 590 68 593 78
rect 617 75 621 78
rect 583 65 593 68
rect 609 67 613 71
rect 647 71 660 75
rect 667 68 670 93
rect 729 93 739 96
rect 701 85 728 89
rect 736 82 739 93
rect 755 95 759 99
rect 763 82 767 87
rect 776 82 780 109
rect 807 93 816 96
rect 790 85 806 89
rect 678 78 714 82
rect 736 78 756 82
rect 763 78 792 82
rect 697 71 728 75
rect 603 64 627 67
rect 661 65 670 68
rect 736 68 739 78
rect 763 75 767 78
rect 729 65 739 68
rect 755 67 759 71
rect 793 71 806 75
rect 813 68 816 93
rect 835 95 839 116
rect 865 112 869 116
rect 907 102 911 116
rect 943 112 947 116
rect 1011 112 1015 116
rect 901 99 925 102
rect 881 93 891 96
rect 833 78 836 82
rect 843 75 847 87
rect 854 85 880 89
rect 888 82 891 93
rect 907 95 911 99
rect 915 82 919 87
rect 928 82 932 109
rect 1053 102 1057 116
rect 1089 112 1093 116
rect 1047 99 1071 102
rect 959 93 968 96
rect 942 85 958 89
rect 854 78 866 82
rect 888 78 908 82
rect 915 78 944 82
rect 847 71 880 75
rect 567 53 571 57
rect 609 53 613 64
rect 749 64 773 67
rect 807 65 816 68
rect 645 53 649 57
rect 713 53 717 57
rect 755 53 759 64
rect 791 53 795 57
rect 835 53 839 71
rect 888 68 891 78
rect 915 75 919 78
rect 881 65 891 68
rect 907 67 911 71
rect 945 71 958 75
rect 965 68 968 93
rect 1027 93 1037 96
rect 999 85 1026 89
rect 1034 82 1037 93
rect 1053 95 1057 99
rect 1061 82 1065 87
rect 1074 82 1078 109
rect 1105 93 1114 96
rect 1088 85 1104 89
rect 976 78 1012 82
rect 1034 78 1054 82
rect 1061 78 1090 82
rect 995 71 1026 75
rect 901 64 925 67
rect 959 65 968 68
rect 1034 68 1037 78
rect 1061 75 1065 78
rect 1027 65 1037 68
rect 1053 67 1057 71
rect 1091 71 1104 75
rect 1111 68 1114 93
rect 865 53 869 57
rect 907 53 911 64
rect 1047 64 1071 67
rect 1105 65 1114 68
rect 943 53 947 57
rect 1011 53 1015 57
rect 1053 53 1057 64
rect 1089 53 1093 57
rect 1948 55 1952 116
rect -65 50 1131 53
rect -77 15 1131 18
rect -61 -6 -57 15
rect -29 11 -25 15
rect 13 -2 17 15
rect 49 11 53 15
rect 117 11 121 15
rect -13 -8 -3 -5
rect -63 -23 -60 -19
rect -53 -26 -49 -14
rect -40 -16 -14 -12
rect -6 -19 -3 -8
rect 34 -19 38 8
rect 159 1 163 15
rect 195 11 199 15
rect 153 -2 177 1
rect 65 -8 74 -5
rect 48 -16 64 -12
rect -40 -23 -28 -19
rect -6 -23 10 -19
rect 30 -23 50 -19
rect -49 -30 -14 -26
rect -61 -48 -57 -30
rect -6 -33 -3 -23
rect 51 -30 64 -26
rect 71 -33 74 -8
rect 133 -8 143 -5
rect 105 -16 132 -12
rect 140 -19 143 -8
rect 159 -6 163 -2
rect 167 -19 171 -14
rect 180 -19 184 8
rect 238 9 242 15
rect 269 11 273 15
rect 211 -8 220 -5
rect 236 -8 239 -4
rect 194 -16 210 -12
rect 82 -23 118 -19
rect 140 -23 160 -19
rect 167 -23 196 -19
rect 101 -30 132 -26
rect -13 -36 -3 -33
rect -29 -48 -25 -44
rect 13 -48 17 -33
rect 65 -36 74 -33
rect 140 -33 143 -23
rect 167 -26 171 -23
rect 133 -36 143 -33
rect 159 -34 163 -30
rect 197 -30 210 -26
rect 217 -33 220 -8
rect 246 -11 250 1
rect 311 1 315 15
rect 347 11 351 15
rect 415 11 419 15
rect 305 -2 329 1
rect 153 -37 177 -34
rect 211 -36 220 -33
rect 49 -48 53 -44
rect 117 -48 121 -44
rect 159 -48 163 -37
rect 195 -48 199 -44
rect 238 -48 242 -15
rect 285 -8 295 -5
rect 246 -26 250 -15
rect 258 -16 284 -12
rect 292 -19 295 -8
rect 311 -6 315 -2
rect 319 -19 323 -14
rect 332 -19 336 8
rect 457 1 461 15
rect 493 11 497 15
rect 451 -2 475 1
rect 363 -8 372 -5
rect 346 -16 362 -12
rect 258 -23 270 -19
rect 292 -23 312 -19
rect 319 -23 348 -19
rect 246 -30 284 -26
rect 292 -33 295 -23
rect 319 -26 323 -23
rect 285 -36 295 -33
rect 311 -34 315 -30
rect 349 -30 362 -26
rect 369 -33 372 -8
rect 431 -8 441 -5
rect 403 -16 430 -12
rect 438 -19 441 -8
rect 457 -6 461 -2
rect 465 -19 469 -14
rect 478 -19 482 8
rect 536 9 540 15
rect 567 11 571 15
rect 509 -8 518 -5
rect 534 -8 537 -4
rect 492 -16 508 -12
rect 380 -23 416 -19
rect 438 -23 458 -19
rect 465 -23 494 -19
rect 399 -30 430 -26
rect 305 -37 329 -34
rect 363 -36 372 -33
rect 438 -33 441 -23
rect 465 -26 469 -23
rect 431 -36 441 -33
rect 457 -34 461 -30
rect 495 -30 508 -26
rect 515 -33 518 -8
rect 544 -11 548 1
rect 609 1 613 15
rect 645 11 649 15
rect 713 11 717 15
rect 603 -2 627 1
rect 269 -48 273 -44
rect 311 -48 315 -37
rect 451 -37 475 -34
rect 509 -36 518 -33
rect 347 -48 351 -44
rect 415 -48 419 -44
rect 457 -48 461 -37
rect 493 -48 497 -44
rect 536 -48 540 -15
rect 583 -8 593 -5
rect 544 -26 548 -15
rect 556 -16 582 -12
rect 590 -19 593 -8
rect 609 -6 613 -2
rect 617 -19 621 -14
rect 630 -19 634 8
rect 755 1 759 15
rect 791 11 795 15
rect 749 -2 773 1
rect 661 -8 670 -5
rect 644 -16 660 -12
rect 556 -23 568 -19
rect 590 -23 610 -19
rect 617 -23 646 -19
rect 544 -30 582 -26
rect 590 -33 593 -23
rect 617 -26 621 -23
rect 583 -36 593 -33
rect 609 -34 613 -30
rect 647 -30 660 -26
rect 667 -33 670 -8
rect 729 -8 739 -5
rect 701 -16 728 -12
rect 736 -19 739 -8
rect 755 -6 759 -2
rect 763 -19 767 -14
rect 776 -19 780 8
rect 834 9 838 15
rect 865 11 869 15
rect 807 -8 816 -5
rect 832 -8 835 -4
rect 790 -16 806 -12
rect 678 -23 714 -19
rect 736 -23 756 -19
rect 763 -23 792 -19
rect 697 -30 728 -26
rect 603 -37 627 -34
rect 661 -36 670 -33
rect 736 -33 739 -23
rect 763 -26 767 -23
rect 729 -36 739 -33
rect 755 -34 759 -30
rect 793 -30 806 -26
rect 813 -33 816 -8
rect 842 -11 846 1
rect 907 1 911 15
rect 943 11 947 15
rect 1011 11 1015 15
rect 901 -2 925 1
rect 567 -48 571 -44
rect 609 -48 613 -37
rect 749 -37 773 -34
rect 807 -36 816 -33
rect 645 -48 649 -44
rect 713 -48 717 -44
rect 755 -48 759 -37
rect 791 -48 795 -44
rect 834 -48 838 -15
rect 881 -8 891 -5
rect 842 -26 846 -15
rect 854 -16 880 -12
rect 888 -19 891 -8
rect 907 -6 911 -2
rect 915 -19 919 -14
rect 928 -19 932 8
rect 1053 1 1057 15
rect 1089 11 1093 15
rect 1047 -2 1071 1
rect 959 -8 968 -5
rect 942 -16 958 -12
rect 854 -23 866 -19
rect 888 -23 908 -19
rect 915 -23 944 -19
rect 842 -30 880 -26
rect 888 -33 891 -23
rect 915 -26 919 -23
rect 881 -36 891 -33
rect 907 -34 911 -30
rect 945 -30 958 -26
rect 965 -33 968 -8
rect 1027 -8 1037 -5
rect 999 -16 1026 -12
rect 1034 -19 1037 -8
rect 1053 -6 1057 -2
rect 1061 -19 1065 -14
rect 1074 -19 1078 8
rect 1105 -8 1114 -5
rect 1088 -16 1104 -12
rect 976 -23 1012 -19
rect 1034 -23 1054 -19
rect 1061 -23 1090 -19
rect 995 -30 1026 -26
rect 901 -37 925 -34
rect 959 -36 968 -33
rect 1034 -33 1037 -23
rect 1061 -26 1065 -23
rect 1027 -36 1037 -33
rect 1053 -34 1057 -30
rect 1091 -30 1104 -26
rect 1111 -33 1114 -8
rect 865 -48 869 -44
rect 907 -48 911 -37
rect 1047 -37 1071 -34
rect 1105 -36 1114 -33
rect 943 -48 947 -44
rect 1011 -48 1015 -44
rect 1053 -48 1057 -37
rect 1089 -48 1093 -44
rect 1948 -48 1952 50
rect 1956 18 1960 116
rect 1972 95 1976 116
rect 2004 112 2008 116
rect 2046 102 2050 116
rect 2082 112 2086 116
rect 2150 112 2154 116
rect 2040 99 2064 102
rect 2020 93 2030 96
rect 1969 78 1973 82
rect 1980 75 1984 87
rect 1993 85 2019 89
rect 2027 82 2030 93
rect 2046 95 2050 99
rect 2054 82 2058 87
rect 2067 82 2071 109
rect 2192 102 2196 116
rect 2228 112 2232 116
rect 2186 99 2210 102
rect 2098 93 2107 96
rect 2081 85 2097 89
rect 1993 78 2005 82
rect 2027 78 2047 82
rect 2054 78 2083 82
rect 1984 71 2019 75
rect 1972 54 1976 71
rect 2027 68 2030 78
rect 2054 75 2058 78
rect 2020 65 2030 68
rect 2046 67 2050 71
rect 2084 71 2097 75
rect 2104 68 2107 93
rect 2166 93 2176 96
rect 2138 85 2165 89
rect 2173 82 2176 93
rect 2192 95 2196 99
rect 2200 82 2204 87
rect 2213 82 2217 109
rect 2244 93 2253 96
rect 2227 85 2243 89
rect 2115 78 2151 82
rect 2173 78 2193 82
rect 2200 78 2229 82
rect 2134 71 2165 75
rect 1968 53 1976 54
rect 2040 64 2064 67
rect 2098 65 2107 68
rect 2173 68 2176 78
rect 2200 75 2204 78
rect 2166 65 2176 68
rect 2192 67 2196 71
rect 2230 71 2243 75
rect 2250 68 2253 93
rect 2272 95 2276 116
rect 2302 112 2306 116
rect 2344 102 2348 116
rect 2380 112 2384 116
rect 2448 112 2452 116
rect 2338 99 2362 102
rect 2318 93 2328 96
rect 2270 78 2273 82
rect 2280 75 2284 87
rect 2291 85 2317 89
rect 2325 82 2328 93
rect 2344 95 2348 99
rect 2352 82 2356 87
rect 2365 82 2369 109
rect 2490 102 2494 116
rect 2526 112 2530 116
rect 2484 99 2508 102
rect 2396 93 2405 96
rect 2379 85 2395 89
rect 2291 78 2303 82
rect 2325 78 2345 82
rect 2352 78 2381 82
rect 2284 71 2317 75
rect 2004 53 2008 57
rect 2046 53 2050 64
rect 2186 64 2210 67
rect 2244 65 2253 68
rect 2082 53 2086 57
rect 2150 53 2154 57
rect 2192 53 2196 64
rect 2228 53 2232 57
rect 2272 53 2276 71
rect 2325 68 2328 78
rect 2352 75 2356 78
rect 2318 65 2328 68
rect 2344 67 2348 71
rect 2382 71 2395 75
rect 2402 68 2405 93
rect 2464 93 2474 96
rect 2436 85 2463 89
rect 2471 82 2474 93
rect 2490 95 2494 99
rect 2498 82 2502 87
rect 2511 82 2515 109
rect 2542 93 2551 96
rect 2525 85 2541 89
rect 2413 78 2449 82
rect 2471 78 2491 82
rect 2498 78 2527 82
rect 2432 71 2463 75
rect 2338 64 2362 67
rect 2396 65 2405 68
rect 2471 68 2474 78
rect 2498 75 2502 78
rect 2464 65 2474 68
rect 2490 67 2494 71
rect 2528 71 2541 75
rect 2548 68 2551 93
rect 2302 53 2306 57
rect 2344 53 2348 64
rect 2484 64 2508 67
rect 2542 65 2551 68
rect 2380 53 2384 57
rect 2448 53 2452 57
rect 2490 53 2494 64
rect 2526 53 2530 57
rect 1968 50 2577 53
rect 1956 15 2577 18
rect 1972 -6 1976 15
rect 2004 11 2008 15
rect 2046 1 2050 15
rect 2082 11 2086 15
rect 2150 11 2154 15
rect 2040 -2 2064 1
rect 2020 -8 2030 -5
rect 1970 -23 1973 -19
rect 1980 -26 1984 -14
rect 1993 -16 2019 -12
rect 2027 -19 2030 -8
rect 2046 -6 2050 -2
rect 2054 -19 2058 -14
rect 2067 -19 2071 8
rect 2192 1 2196 15
rect 2228 11 2232 15
rect 2186 -2 2210 1
rect 2098 -8 2107 -5
rect 2081 -16 2097 -12
rect 1993 -23 2005 -19
rect 2027 -23 2047 -19
rect 2054 -23 2083 -19
rect 1984 -30 2019 -26
rect 1972 -48 1976 -30
rect 2027 -33 2030 -23
rect 2054 -26 2058 -23
rect 2020 -36 2030 -33
rect 2046 -34 2050 -30
rect 2084 -30 2097 -26
rect 2104 -33 2107 -8
rect 2166 -8 2176 -5
rect 2138 -16 2165 -12
rect 2173 -19 2176 -8
rect 2192 -6 2196 -2
rect 2200 -19 2204 -14
rect 2213 -19 2217 8
rect 2271 9 2275 15
rect 2302 11 2306 15
rect 2244 -8 2253 -5
rect 2269 -8 2272 -4
rect 2227 -16 2243 -12
rect 2115 -23 2151 -19
rect 2173 -23 2193 -19
rect 2200 -23 2229 -19
rect 2134 -30 2165 -26
rect 2040 -37 2064 -34
rect 2098 -36 2107 -33
rect 2173 -33 2176 -23
rect 2200 -26 2204 -23
rect 2166 -36 2176 -33
rect 2192 -34 2196 -30
rect 2230 -30 2243 -26
rect 2250 -33 2253 -8
rect 2279 -11 2283 1
rect 2344 1 2348 15
rect 2380 11 2384 15
rect 2448 11 2452 15
rect 2338 -2 2362 1
rect 2004 -48 2008 -44
rect 2046 -48 2050 -37
rect 2186 -37 2210 -34
rect 2244 -36 2253 -33
rect 2082 -48 2086 -44
rect 2150 -48 2154 -44
rect 2192 -48 2196 -37
rect 2228 -48 2232 -44
rect 2271 -48 2275 -15
rect 2318 -8 2328 -5
rect 2279 -26 2283 -15
rect 2291 -16 2317 -12
rect 2325 -19 2328 -8
rect 2344 -6 2348 -2
rect 2352 -19 2356 -14
rect 2365 -19 2369 8
rect 2490 1 2494 15
rect 2526 11 2530 15
rect 2484 -2 2508 1
rect 2396 -8 2405 -5
rect 2379 -16 2395 -12
rect 2291 -23 2303 -19
rect 2325 -23 2345 -19
rect 2352 -23 2381 -19
rect 2279 -30 2317 -26
rect 2325 -33 2328 -23
rect 2352 -26 2356 -23
rect 2318 -36 2328 -33
rect 2344 -34 2348 -30
rect 2382 -30 2395 -26
rect 2402 -33 2405 -8
rect 2464 -8 2474 -5
rect 2436 -16 2463 -12
rect 2471 -19 2474 -8
rect 2490 -6 2494 -2
rect 2498 -19 2502 -14
rect 2511 -19 2515 8
rect 2542 -8 2551 -5
rect 2525 -16 2541 -12
rect 2413 -23 2449 -19
rect 2471 -23 2491 -19
rect 2498 -23 2527 -19
rect 2432 -30 2463 -26
rect 2338 -37 2362 -34
rect 2396 -36 2405 -33
rect 2471 -33 2474 -23
rect 2498 -26 2502 -23
rect 2464 -36 2474 -33
rect 2490 -34 2494 -30
rect 2528 -30 2541 -26
rect 2548 -33 2551 -8
rect 2302 -48 2306 -44
rect 2344 -48 2348 -37
rect 2484 -37 2508 -34
rect 2542 -36 2551 -33
rect 2380 -48 2384 -44
rect 2448 -48 2452 -44
rect 2490 -48 2494 -37
rect 2526 -48 2530 -44
rect -85 -51 2577 -48
rect 2565 -62 2577 -58
rect 1128 -71 1131 -67
rect 2267 -71 2577 -67
rect 830 -79 1131 -75
rect 532 -87 1131 -83
rect 234 -95 1131 -91
<< m2contact >>
rect 1959 190 1964 195
rect 1989 186 1994 191
rect 2064 201 2069 206
rect 2029 170 2034 175
rect 2072 167 2077 172
rect 2135 186 2140 191
rect 2103 175 2108 180
rect 2210 201 2215 206
rect 2122 167 2127 172
rect 2100 162 2105 167
rect 2175 170 2180 175
rect 2218 167 2223 172
rect 2255 170 2260 175
rect 2246 162 2251 167
rect -85 50 -80 55
rect -37 89 -32 94
rect -69 78 -64 83
rect 38 104 43 109
rect -70 50 -65 55
rect 3 73 8 78
rect 46 70 51 75
rect 109 89 114 94
rect 77 78 82 83
rect 96 70 101 75
rect 74 65 79 70
rect 149 73 154 78
rect 192 70 197 75
rect 261 89 266 94
rect 232 78 237 83
rect 336 104 341 109
rect 220 65 225 70
rect 301 73 306 78
rect 344 70 349 75
rect 407 89 412 94
rect 375 78 380 83
rect 394 70 399 75
rect 372 65 377 70
rect 447 73 452 78
rect 490 70 495 75
rect 559 89 564 94
rect 530 78 535 83
rect 634 104 639 109
rect 518 65 523 70
rect 599 73 604 78
rect 642 70 647 75
rect 705 89 710 94
rect 673 78 678 83
rect 692 70 697 75
rect 670 65 675 70
rect 745 73 750 78
rect 788 70 793 75
rect 857 89 862 94
rect 828 78 833 83
rect 932 104 937 109
rect 816 65 821 70
rect 897 73 902 78
rect 940 70 945 75
rect 1003 89 1008 94
rect 971 78 976 83
rect 990 70 995 75
rect 968 65 973 70
rect 1043 73 1048 78
rect 1086 70 1091 75
rect 1114 65 1119 70
rect 1948 50 1953 55
rect -37 -12 -32 -7
rect -68 -23 -63 -18
rect 38 3 43 8
rect 3 -28 8 -23
rect 46 -31 51 -26
rect 109 -12 114 -7
rect 77 -23 82 -18
rect 184 3 189 8
rect 231 -8 236 -3
rect 96 -31 101 -26
rect 74 -36 79 -31
rect 149 -28 154 -23
rect 192 -31 197 -26
rect 220 -36 225 -31
rect 261 -12 266 -7
rect 336 3 341 8
rect 301 -28 306 -23
rect 344 -31 349 -26
rect 407 -12 412 -7
rect 375 -23 380 -18
rect 482 3 487 8
rect 529 -8 534 -3
rect 394 -31 399 -26
rect 372 -36 377 -31
rect 447 -28 452 -23
rect 490 -31 495 -26
rect 518 -36 523 -31
rect 559 -12 564 -7
rect 634 3 639 8
rect 599 -28 604 -23
rect 642 -31 647 -26
rect 705 -12 710 -7
rect 673 -23 678 -18
rect 780 3 785 8
rect 827 -8 832 -3
rect 692 -31 697 -26
rect 670 -36 675 -31
rect 745 -28 750 -23
rect 788 -31 793 -26
rect 816 -36 821 -31
rect 857 -12 862 -7
rect 932 3 937 8
rect 897 -28 902 -23
rect 940 -31 945 -26
rect 1003 -12 1008 -7
rect 971 -23 976 -18
rect 1078 3 1083 8
rect 990 -31 995 -26
rect 968 -36 973 -31
rect 1043 -28 1048 -23
rect 1086 -31 1091 -26
rect 1114 -36 1119 -31
rect 1996 89 2001 94
rect 1964 78 1969 83
rect 2071 104 2076 109
rect 1963 50 1968 55
rect 2036 73 2041 78
rect 2079 70 2084 75
rect 2142 89 2147 94
rect 2110 78 2115 83
rect 2129 70 2134 75
rect 2107 65 2112 70
rect 2182 73 2187 78
rect 2225 70 2230 75
rect 2294 89 2299 94
rect 2265 78 2270 83
rect 2369 104 2374 109
rect 2253 65 2258 70
rect 2334 73 2339 78
rect 2377 70 2382 75
rect 2440 89 2445 94
rect 2408 78 2413 83
rect 2427 70 2432 75
rect 2405 65 2410 70
rect 2480 73 2485 78
rect 2523 70 2528 75
rect 2551 65 2556 70
rect 1996 -12 2001 -7
rect 1965 -23 1970 -18
rect 2071 3 2076 8
rect 2036 -28 2041 -23
rect 2079 -31 2084 -26
rect 2142 -12 2147 -7
rect 2110 -23 2115 -18
rect 2217 3 2222 8
rect 2264 -8 2269 -3
rect 2129 -31 2134 -26
rect 2107 -36 2112 -31
rect 2182 -28 2187 -23
rect 2225 -31 2230 -26
rect 2253 -36 2258 -31
rect 2294 -12 2299 -7
rect 2369 3 2374 8
rect 2334 -28 2339 -23
rect 2377 -31 2382 -26
rect 2440 -12 2445 -7
rect 2408 -23 2413 -18
rect 2515 3 2520 8
rect 2427 -31 2432 -26
rect 2405 -36 2410 -31
rect 2480 -28 2485 -23
rect 2523 -31 2528 -26
rect 2551 -36 2556 -31
rect 2560 -63 2565 -58
rect 1123 -71 1128 -66
rect 2262 -71 2267 -66
rect 825 -79 830 -74
rect 527 -87 532 -82
rect 229 -95 234 -90
<< metal2 >>
rect 2056 226 2122 230
rect 2056 222 2060 226
rect 1959 218 2060 222
rect 1959 195 1963 218
rect 1989 191 1993 218
rect 2056 172 2060 218
rect 2065 218 2107 222
rect 2065 206 2069 218
rect 2103 180 2107 218
rect 2029 145 2033 170
rect 2056 168 2072 172
rect 2118 168 2122 226
rect 2135 218 2206 222
rect 2135 191 2139 218
rect 2202 172 2206 218
rect 2211 218 2253 222
rect 2211 206 2215 218
rect 2249 175 2253 218
rect 2100 145 2104 162
rect 2029 141 2104 145
rect 2175 145 2179 170
rect 2202 168 2218 172
rect 2249 171 2255 175
rect 2246 145 2250 162
rect 2175 141 2250 145
rect 30 129 96 133
rect 30 125 34 129
rect -69 121 34 125
rect -69 83 -65 121
rect -37 94 -33 121
rect 30 75 34 121
rect 39 121 81 125
rect 39 109 43 121
rect 77 83 81 121
rect -80 50 -70 54
rect 3 48 7 73
rect 30 71 46 75
rect 92 71 96 129
rect 328 129 394 133
rect 328 125 332 129
rect 109 121 180 125
rect 109 94 113 121
rect 176 75 180 121
rect 261 121 332 125
rect 261 106 265 121
rect 232 102 265 106
rect 232 83 236 102
rect 261 94 265 102
rect 74 48 78 65
rect 3 44 78 48
rect 149 48 153 73
rect 176 71 192 75
rect 328 75 332 121
rect 337 121 379 125
rect 337 109 341 121
rect 375 83 379 121
rect 220 48 224 65
rect 149 44 224 48
rect 301 48 305 73
rect 328 71 344 75
rect 390 71 394 129
rect 626 129 692 133
rect 626 125 630 129
rect 407 121 478 125
rect 407 94 411 121
rect 474 75 478 121
rect 559 121 630 125
rect 559 106 563 121
rect 530 102 563 106
rect 530 83 534 102
rect 559 94 563 102
rect 372 48 376 65
rect 301 44 376 48
rect 447 48 451 73
rect 474 71 490 75
rect 626 75 630 121
rect 635 121 677 125
rect 635 109 639 121
rect 673 83 677 121
rect 518 48 522 65
rect 447 44 522 48
rect 599 48 603 73
rect 626 71 642 75
rect 688 71 692 129
rect 924 129 990 133
rect 924 125 928 129
rect 705 121 776 125
rect 705 94 709 121
rect 772 75 776 121
rect 857 121 928 125
rect 857 106 861 121
rect 828 102 861 106
rect 828 83 832 102
rect 857 94 861 102
rect 670 48 674 65
rect 599 44 674 48
rect 745 48 749 73
rect 772 71 788 75
rect 924 75 928 121
rect 933 121 975 125
rect 933 109 937 121
rect 971 83 975 121
rect 816 48 820 65
rect 745 44 820 48
rect 897 48 901 73
rect 924 71 940 75
rect 986 71 990 129
rect 2063 129 2129 133
rect 2063 125 2067 129
rect 1003 121 1074 125
rect 1003 94 1007 121
rect 1070 75 1074 121
rect 1964 121 2067 125
rect 1964 83 1968 121
rect 1996 94 2000 121
rect 968 48 972 65
rect 897 44 972 48
rect 1043 48 1047 73
rect 1070 71 1086 75
rect 2063 75 2067 121
rect 2072 121 2114 125
rect 2072 109 2076 121
rect 2110 83 2114 121
rect 1114 48 1118 65
rect 1953 50 1963 54
rect 1043 44 1118 48
rect 2036 48 2040 73
rect 2063 71 2079 75
rect 2125 71 2129 129
rect 2361 129 2427 133
rect 2361 125 2365 129
rect 2142 121 2213 125
rect 2142 94 2146 121
rect 2209 75 2213 121
rect 2294 121 2365 125
rect 2294 106 2298 121
rect 2265 102 2298 106
rect 2265 83 2269 102
rect 2294 94 2298 102
rect 2107 48 2111 65
rect 2036 44 2111 48
rect 2182 48 2186 73
rect 2209 71 2225 75
rect 2361 75 2365 121
rect 2370 121 2412 125
rect 2370 109 2374 121
rect 2408 83 2412 121
rect 2253 48 2257 65
rect 2182 44 2257 48
rect 2334 48 2338 73
rect 2361 71 2377 75
rect 2423 71 2427 129
rect 2440 121 2511 125
rect 2440 94 2444 121
rect 2507 75 2511 121
rect 2405 48 2409 65
rect 2334 44 2409 48
rect 2480 48 2484 73
rect 2507 71 2523 75
rect 2551 48 2555 65
rect 2480 44 2555 48
rect 30 28 96 32
rect 30 24 34 28
rect -68 20 34 24
rect -68 -18 -64 20
rect -37 -7 -33 20
rect 30 -26 34 20
rect 39 20 81 24
rect 39 8 43 20
rect 77 -18 81 20
rect 3 -53 7 -28
rect 30 -30 46 -26
rect 92 -30 96 28
rect 328 28 394 32
rect 328 24 332 28
rect 109 20 180 24
rect 109 -7 113 20
rect 176 -26 180 20
rect 185 20 227 24
rect 185 8 189 20
rect 223 -23 227 20
rect 231 20 332 24
rect 231 -3 235 20
rect 261 -7 265 20
rect 74 -53 78 -36
rect 3 -57 78 -53
rect 149 -53 153 -28
rect 176 -30 192 -26
rect 223 -27 233 -23
rect 220 -53 224 -36
rect 149 -57 224 -53
rect 229 -90 233 -27
rect 328 -26 332 20
rect 337 20 379 24
rect 337 8 341 20
rect 375 -18 379 20
rect 301 -53 305 -28
rect 328 -30 344 -26
rect 390 -30 394 28
rect 626 28 692 32
rect 626 24 630 28
rect 407 20 478 24
rect 407 -7 411 20
rect 474 -26 478 20
rect 483 20 525 24
rect 483 8 487 20
rect 521 -23 525 20
rect 529 20 630 24
rect 529 -3 533 20
rect 559 -7 563 20
rect 372 -53 376 -36
rect 301 -57 376 -53
rect 447 -53 451 -28
rect 474 -30 490 -26
rect 521 -27 531 -23
rect 518 -53 522 -36
rect 447 -57 522 -53
rect 527 -82 531 -27
rect 626 -26 630 20
rect 635 20 677 24
rect 635 8 639 20
rect 673 -18 677 20
rect 599 -53 603 -28
rect 626 -30 642 -26
rect 688 -30 692 28
rect 924 28 990 32
rect 924 24 928 28
rect 705 20 776 24
rect 705 -7 709 20
rect 772 -26 776 20
rect 781 20 823 24
rect 781 8 785 20
rect 819 -23 823 20
rect 827 20 928 24
rect 827 -3 831 20
rect 857 -7 861 20
rect 670 -53 674 -36
rect 599 -57 674 -53
rect 745 -53 749 -28
rect 772 -30 788 -26
rect 819 -27 829 -23
rect 816 -53 820 -36
rect 745 -57 820 -53
rect 825 -74 829 -27
rect 924 -26 928 20
rect 933 20 975 24
rect 933 8 937 20
rect 971 -18 975 20
rect 897 -53 901 -28
rect 924 -30 940 -26
rect 986 -30 990 28
rect 2063 28 2129 32
rect 2063 24 2067 28
rect 1003 20 1074 24
rect 1003 -7 1007 20
rect 1070 -26 1074 20
rect 1079 20 1121 24
rect 1079 8 1083 20
rect 1117 -23 1121 20
rect 1965 20 2067 24
rect 1965 -18 1969 20
rect 1996 -7 2000 20
rect 968 -53 972 -36
rect 897 -57 972 -53
rect 1043 -53 1047 -28
rect 1070 -30 1086 -26
rect 1117 -27 1127 -23
rect 1114 -53 1118 -36
rect 1043 -57 1118 -53
rect 1123 -66 1127 -27
rect 2063 -26 2067 20
rect 2072 20 2114 24
rect 2072 8 2076 20
rect 2110 -18 2114 20
rect 2036 -53 2040 -28
rect 2063 -30 2079 -26
rect 2125 -30 2129 28
rect 2361 28 2427 32
rect 2361 24 2365 28
rect 2142 20 2213 24
rect 2142 -7 2146 20
rect 2209 -26 2213 20
rect 2218 20 2260 24
rect 2218 8 2222 20
rect 2256 -23 2260 20
rect 2264 20 2365 24
rect 2264 -3 2268 20
rect 2294 -7 2298 20
rect 2107 -53 2111 -36
rect 2036 -57 2111 -53
rect 2182 -53 2186 -28
rect 2209 -30 2225 -26
rect 2256 -27 2266 -23
rect 2253 -53 2257 -36
rect 2182 -57 2257 -53
rect 2262 -66 2266 -27
rect 2361 -26 2365 20
rect 2370 20 2412 24
rect 2370 8 2374 20
rect 2408 -18 2412 20
rect 2334 -53 2338 -28
rect 2361 -30 2377 -26
rect 2423 -30 2427 28
rect 2440 20 2511 24
rect 2440 -7 2444 20
rect 2507 -26 2511 20
rect 2516 20 2558 24
rect 2516 8 2520 20
rect 2554 -23 2558 20
rect 2405 -53 2409 -36
rect 2334 -57 2409 -53
rect 2480 -53 2484 -28
rect 2507 -30 2523 -26
rect 2554 -27 2564 -23
rect 2551 -53 2555 -36
rect 2480 -57 2555 -53
rect 2560 -58 2564 -27
<< m123contact >>
rect 2069 182 2074 187
rect 229 160 234 165
rect 1989 163 1994 168
rect 527 152 532 157
rect 825 144 830 149
rect 2126 182 2131 187
rect 2215 182 2220 187
rect 2135 163 2140 168
rect 1123 137 1128 142
rect 2262 136 2267 141
rect 43 85 48 90
rect -37 66 -32 71
rect 100 85 105 90
rect 184 104 189 109
rect 189 85 194 90
rect 109 66 114 71
rect 341 85 346 90
rect 261 66 266 71
rect 398 85 403 90
rect 482 104 487 109
rect 487 85 492 90
rect 407 66 412 71
rect 639 85 644 90
rect 559 66 564 71
rect 696 85 701 90
rect 780 104 785 109
rect 785 85 790 90
rect 705 66 710 71
rect 937 85 942 90
rect 857 66 862 71
rect 994 85 999 90
rect 1078 104 1083 109
rect 1083 85 1088 90
rect 1003 66 1008 71
rect 2076 85 2081 90
rect 1996 66 2001 71
rect 2133 85 2138 90
rect 2217 104 2222 109
rect 2222 85 2227 90
rect 2142 66 2147 71
rect 2374 85 2379 90
rect 2294 66 2299 71
rect 2516 122 2521 127
rect 2431 85 2436 90
rect 2515 104 2520 109
rect 2520 85 2525 90
rect 2440 66 2445 71
rect 43 -16 48 -11
rect -37 -35 -32 -30
rect 100 -16 105 -11
rect 189 -16 194 -11
rect 109 -35 114 -30
rect 341 -16 346 -11
rect 261 -35 266 -30
rect 398 -16 403 -11
rect 487 -16 492 -11
rect 407 -35 412 -30
rect 639 -16 644 -11
rect 559 -35 564 -30
rect 696 -16 701 -11
rect 785 -16 790 -11
rect 705 -35 710 -30
rect 937 -16 942 -11
rect 857 -35 862 -30
rect 994 -16 999 -11
rect 1083 -16 1088 -11
rect 1003 -35 1008 -30
rect 2076 -16 2081 -11
rect 1996 -35 2001 -30
rect 2133 -16 2138 -11
rect 2222 -16 2227 -11
rect 2142 -35 2147 -30
rect 2374 -16 2379 -11
rect 2294 -35 2299 -30
rect 2431 -16 2436 -11
rect 2520 -16 2525 -11
rect 2440 -35 2445 -30
<< metal3 >>
rect 229 125 233 160
rect 527 125 531 152
rect 825 125 829 144
rect 1989 139 1993 163
rect 2065 158 2069 187
rect 2112 182 2126 186
rect 2021 154 2069 158
rect 2021 139 2025 154
rect 2112 139 2116 182
rect 2135 146 2139 163
rect 2211 158 2215 187
rect 2167 154 2215 158
rect 2167 146 2171 154
rect 2135 143 2171 146
rect 1123 125 1127 137
rect 1989 135 2116 139
rect 2262 125 2266 136
rect 185 121 233 125
rect 483 121 531 125
rect 781 121 829 125
rect 1079 121 1127 125
rect 2218 121 2266 125
rect 185 109 189 121
rect 483 109 487 121
rect 781 109 785 121
rect 1079 109 1083 121
rect 2218 109 2222 121
rect 2516 109 2520 122
rect -37 48 -33 66
rect 39 61 43 90
rect 86 85 100 89
rect -5 57 43 61
rect -5 48 -1 57
rect -37 44 -1 48
rect -5 42 -1 44
rect 86 42 90 85
rect 109 49 113 66
rect 185 61 189 90
rect 141 57 189 61
rect 141 49 145 57
rect 109 46 145 49
rect -5 38 90 42
rect 261 42 265 66
rect 337 61 341 90
rect 384 85 398 89
rect 293 57 341 61
rect 293 42 297 57
rect 384 42 388 85
rect 407 49 411 66
rect 483 61 487 90
rect 439 57 487 61
rect 439 49 443 57
rect 407 46 443 49
rect 261 38 388 42
rect 559 42 563 66
rect 635 61 639 90
rect 682 85 696 89
rect 591 57 639 61
rect 591 42 595 57
rect 682 42 686 85
rect 705 49 709 66
rect 781 61 785 90
rect 737 57 785 61
rect 737 49 741 57
rect 705 46 741 49
rect 559 38 686 42
rect 857 42 861 66
rect 933 61 937 90
rect 980 85 994 89
rect 889 57 937 61
rect 889 42 893 57
rect 980 42 984 85
rect 1003 49 1007 66
rect 1079 61 1083 90
rect 1035 57 1083 61
rect 1035 49 1039 57
rect 1003 46 1039 49
rect 1996 48 2000 66
rect 2072 61 2076 90
rect 2119 85 2133 89
rect 2028 57 2076 61
rect 2028 48 2032 57
rect 1996 44 2032 48
rect 857 38 984 42
rect 2028 42 2032 44
rect 2119 42 2123 85
rect 2142 49 2146 66
rect 2218 61 2222 90
rect 2174 57 2222 61
rect 2174 49 2178 57
rect 2142 46 2178 49
rect 2028 38 2123 42
rect 2294 42 2298 66
rect 2370 61 2374 90
rect 2417 85 2431 89
rect 2326 57 2374 61
rect 2326 42 2330 57
rect 2417 42 2421 85
rect 2440 49 2444 66
rect 2516 61 2520 90
rect 2472 57 2520 61
rect 2472 49 2476 57
rect 2440 46 2476 49
rect 2294 38 2421 42
rect -37 -53 -33 -35
rect 39 -40 43 -11
rect 86 -16 100 -12
rect -5 -44 43 -40
rect -5 -53 -1 -44
rect -37 -57 -1 -53
rect -5 -59 -1 -57
rect 86 -59 90 -16
rect 109 -52 113 -35
rect 185 -40 189 -11
rect 141 -44 189 -40
rect 141 -52 145 -44
rect 109 -55 145 -52
rect -5 -63 90 -59
rect 261 -59 265 -35
rect 337 -40 341 -11
rect 384 -16 398 -12
rect 293 -44 341 -40
rect 293 -59 297 -44
rect 384 -59 388 -16
rect 407 -52 411 -35
rect 483 -40 487 -11
rect 439 -44 487 -40
rect 439 -52 443 -44
rect 407 -55 443 -52
rect 261 -63 388 -59
rect 559 -59 563 -35
rect 635 -40 639 -11
rect 682 -16 696 -12
rect 591 -44 639 -40
rect 591 -59 595 -44
rect 682 -59 686 -16
rect 705 -52 709 -35
rect 781 -40 785 -11
rect 737 -44 785 -40
rect 737 -52 741 -44
rect 705 -55 741 -52
rect 559 -63 686 -59
rect 857 -59 861 -35
rect 933 -40 937 -11
rect 980 -16 994 -12
rect 889 -44 937 -40
rect 889 -59 893 -44
rect 980 -59 984 -16
rect 1003 -52 1007 -35
rect 1079 -40 1083 -11
rect 1035 -44 1083 -40
rect 1035 -52 1039 -44
rect 1003 -55 1039 -52
rect 1996 -53 2000 -35
rect 2072 -40 2076 -11
rect 2119 -16 2133 -12
rect 2028 -44 2076 -40
rect 2028 -53 2032 -44
rect 1996 -57 2032 -53
rect 857 -63 984 -59
rect 2028 -59 2032 -57
rect 2119 -59 2123 -16
rect 2142 -52 2146 -35
rect 2218 -40 2222 -11
rect 2174 -44 2222 -40
rect 2174 -52 2178 -44
rect 2142 -55 2178 -52
rect 2028 -63 2123 -59
rect 2294 -59 2298 -35
rect 2370 -40 2374 -11
rect 2417 -16 2431 -12
rect 2326 -44 2374 -40
rect 2326 -59 2330 -44
rect 2417 -59 2421 -16
rect 2440 -52 2444 -35
rect 2516 -40 2520 -11
rect 2472 -44 2520 -40
rect 2472 -52 2476 -44
rect 2440 -55 2476 -52
rect 2294 -63 2421 -59
use MNSinv  MNSinv_0
timestamp 1618889747
transform 1 0 26 0 1 -17
box -19 -20 5 18
<< labels >>
rlabel metal1 159 101 170 102 5 vdd
rlabel metal1 163 64 167 65 1 gnd
rlabel metal1 13 101 24 102 5 vdd
rlabel metal1 17 64 21 65 1 gnd
rlabel metal1 -38 -22 -35 -21 1 a3_d
rlabel ndcontact -20 -42 -18 -41 1 a302
rlabel pdcontact -20 1 -18 2 1 a301
rlabel metal1 -2 -22 2 -21 1 a303
rlabel metal1 35 -22 37 -21 1 a304
rlabel pdcontact 58 1 60 2 1 a305
rlabel ndcontact 58 -42 60 -41 1 a306
rlabel ndcontact 126 -42 128 -41 1 a308
rlabel pdcontact 126 1 128 2 1 a307
rlabel metal1 144 -22 148 -21 1 a309
rlabel pdcontact 204 1 206 2 1 a310
rlabel ndcontact 204 -42 206 -41 1 a311
rlabel metal1 181 -22 184 -21 1 a3
rlabel ndcontact 204 59 206 60 1 b311
rlabel pdcontact 204 102 206 103 1 b310
rlabel metal1 181 79 184 80 1 b3
rlabel metal1 144 79 148 80 1 b309
rlabel ndcontact 126 59 128 60 1 b308
rlabel pdcontact 126 102 128 103 1 b307
rlabel ndcontact 58 59 60 60 1 b306
rlabel pdcontact 58 102 60 103 1 b305
rlabel metal1 35 79 38 80 1 b304
rlabel metal1 -2 79 2 80 1 b303
rlabel ndcontact -20 59 -18 60 1 b302
rlabel pdcontact -20 102 -18 103 1 b301
rlabel metal1 -37 79 -34 80 1 b3_d
rlabel metal1 457 101 468 102 5 vdd
rlabel metal1 461 64 465 65 1 gnd
rlabel metal1 311 101 322 102 5 vdd
rlabel metal1 315 64 319 65 1 gnd
rlabel metal1 261 -22 264 -21 1 a2_d
rlabel ndcontact 502 -42 504 -41 1 a211
rlabel pdcontact 502 1 504 2 1 a210
rlabel ndcontact 424 -42 426 -41 1 a208
rlabel pdcontact 424 1 426 2 1 a207
rlabel ndcontact 356 -42 358 -41 1 a206
rlabel pdcontact 356 1 358 2 1 a205
rlabel ndcontact 278 -42 280 -41 1 a202
rlabel pdcontact 278 1 280 2 1 a201
rlabel metal1 296 -22 300 -21 1 a203
rlabel metal1 333 -22 336 -21 1 a204
rlabel metal1 442 -22 446 -21 1 a209
rlabel metal1 479 -22 482 -21 1 a2
rlabel metal1 479 79 482 80 1 b2
rlabel metal1 442 79 446 80 1 b209
rlabel metal1 296 79 300 80 1 b203
rlabel metal1 333 79 336 80 1 b204
rlabel metal1 261 79 264 80 1 b2_d
rlabel pdcontact 278 102 280 103 1 b201
rlabel ndcontact 278 59 280 60 1 b202
rlabel pdcontact 356 102 358 103 1 b205
rlabel ndcontact 356 59 358 60 1 b206
rlabel pdcontact 424 102 426 103 1 b207
rlabel ndcontact 424 59 426 60 1 b208
rlabel pdcontact 502 102 504 103 1 b210
rlabel ndcontact 502 59 504 60 1 b211
rlabel metal1 755 101 766 102 5 vdd
rlabel metal1 759 64 763 65 1 gnd
rlabel metal1 609 101 620 102 5 vdd
rlabel metal1 613 64 617 65 1 gnd
rlabel metal1 559 -22 562 -21 1 a1_d
rlabel pdcontact 576 1 578 2 1 a101
rlabel ndcontact 576 -42 578 -41 1 a102
rlabel pdcontact 654 1 656 2 1 a105
rlabel ndcontact 654 -42 656 -41 1 a106
rlabel pdcontact 722 1 724 2 1 a107
rlabel ndcontact 722 -42 724 -41 1 a108
rlabel pdcontact 800 1 802 2 1 a110
rlabel ndcontact 800 -42 802 -41 1 a111
rlabel metal1 777 -22 780 -21 1 a1
rlabel metal1 740 -22 744 -21 1 a109
rlabel metal1 631 -22 634 -21 1 a104
rlabel metal1 594 -22 598 -21 1 a103
rlabel ndcontact 800 59 802 60 1 b111
rlabel pdcontact 800 102 802 103 1 b110
rlabel ndcontact 722 59 724 60 1 b108
rlabel pdcontact 722 102 724 103 1 b107
rlabel ndcontact 654 59 656 60 1 b106
rlabel pdcontact 654 102 656 103 1 b105
rlabel ndcontact 576 59 578 60 1 b102
rlabel pdcontact 576 102 578 103 1 b101
rlabel metal1 559 79 562 80 1 b1_d
rlabel metal1 594 79 598 80 1 b103
rlabel metal1 631 79 634 80 1 b104
rlabel metal1 740 79 744 80 1 b109
rlabel metal1 777 79 780 80 1 b1
rlabel metal1 1053 0 1064 1 5 vdd
rlabel metal1 1057 -37 1061 -36 1 gnd
rlabel pdcontact 874 1 876 2 1 a001
rlabel ndcontact 874 -42 876 -41 1 a002
rlabel metal1 892 -22 896 -21 1 a003
rlabel metal1 929 -22 932 -21 1 a004
rlabel pdcontact 952 1 954 2 1 a005
rlabel ndcontact 952 -42 954 -41 1 a006
rlabel pdcontact 1020 1 1022 2 1 a007
rlabel ndcontact 1020 -42 1022 -41 1 a008
rlabel metal1 1038 -22 1042 -21 1 a009
rlabel pdcontact 1098 1 1100 2 1 a010
rlabel ndcontact 1098 -42 1100 -41 1 a011
rlabel metal1 857 -22 860 -21 1 a0_d
rlabel metal1 1075 -22 1078 -21 1 a0
rlabel metal1 1053 101 1064 102 5 vdd
rlabel metal1 1057 64 1061 65 1 gnd
rlabel metal1 907 101 918 102 5 vdd
rlabel metal1 911 64 915 65 1 gnd
rlabel metal1 1075 79 1078 80 1 b0
rlabel metal1 1038 79 1042 80 1 b009
rlabel metal1 892 79 896 80 1 b003
rlabel metal1 929 79 932 80 1 b004
rlabel metal1 857 79 860 80 1 b0_d
rlabel ndcontact 874 59 876 60 1 b002
rlabel pdcontact 874 102 876 103 1 b001
rlabel ndcontact 952 59 954 60 1 b006
rlabel pdcontact 952 102 954 103 1 b005
rlabel ndcontact 1020 59 1022 60 1 b008
rlabel pdcontact 1020 102 1022 103 1 b007
rlabel ndcontact 1098 59 1100 60 1 b011
rlabel pdcontact 1098 102 1100 103 1 b010
rlabel metal1 -38 -15 -35 -14 1 clka3
rlabel metal1 -38 -29 -35 -28 1 clka3_bar
rlabel metal1 260 -29 262 -28 1 clka2_bar
rlabel metal1 260 -15 262 -14 1 clka2
rlabel metal1 558 -29 560 -28 1 clka1_bar
rlabel metal1 558 -15 560 -14 1 clka1
rlabel metal1 856 -29 858 -28 1 clka0_bar
rlabel metal1 856 -15 858 -14 1 clka0
rlabel metal1 856 72 858 73 1 clkb0_bar
rlabel metal1 856 86 858 87 1 clkb0
rlabel metal1 558 72 560 73 1 clkb1_bar
rlabel metal1 558 86 560 87 1 clkb1
rlabel metal1 260 72 262 73 1 clkb2_bar
rlabel metal1 260 86 262 87 1 clkb2
rlabel metal1 -38 72 -36 73 1 clkb3_bar
rlabel metal1 -38 86 -36 87 1 clkb3
rlabel metal1 2192 0 2203 1 5 vdd
rlabel metal1 2196 -37 2200 -36 1 gnd
rlabel metal1 2192 101 2203 102 5 vdd
rlabel metal1 2196 64 2200 65 1 gnd
rlabel metal1 2046 101 2057 102 5 vdd
rlabel metal1 2050 64 2054 65 1 gnd
rlabel metal1 2490 0 2501 1 5 vdd
rlabel metal1 2494 -37 2498 -36 1 gnd
rlabel metal1 2490 101 2501 102 5 vdd
rlabel metal1 2494 64 2498 65 1 gnd
rlabel metal1 2344 101 2355 102 5 vdd
rlabel metal1 2348 64 2352 65 1 gnd
rlabel metal1 2344 0 2355 1 5 vdd
rlabel metal1 2348 -37 2352 -36 1 gnd
rlabel metal1 2046 0 2057 1 5 vdd
rlabel metal1 2050 -37 2054 -36 1 gnd
rlabel metal1 1995 -15 1998 -14 1 clks2
rlabel metal1 1995 -22 1998 -21 1 s2
rlabel metal1 1995 -29 1998 -28 1 clks2_bar
rlabel pdcontact 2013 1 2015 2 1 s201
rlabel ndcontact 2013 -42 2015 -41 1 s202
rlabel metal1 2068 -22 2070 -21 1 s204
rlabel pdcontact 2091 1 2093 2 1 s205
rlabel ndcontact 2091 -42 2093 -41 1 s206
rlabel pdcontact 2159 1 2161 2 1 s207
rlabel ndcontact 2159 -42 2161 -41 1 s208
rlabel ndcontact 2237 -42 2239 -41 1 s211
rlabel pdcontact 2237 1 2239 2 1 s210
rlabel metal1 2214 -22 2217 -21 1 s2_q
rlabel metal1 2177 -22 2181 -21 1 s209
rlabel metal1 2031 -22 2035 -21 1 s203
rlabel metal1 2293 -29 2295 -28 1 clks0_bar
rlabel metal1 2293 -15 2295 -14 1 clks0
rlabel metal1 2294 -22 2297 -21 1 s0
rlabel ndcontact 2311 -42 2313 -41 1 s002
rlabel pdcontact 2311 1 2313 2 1 s001
rlabel ndcontact 2389 -42 2391 -41 1 s006
rlabel pdcontact 2389 1 2391 2 1 s005
rlabel ndcontact 2457 -42 2459 -41 1 s008
rlabel pdcontact 2457 1 2459 2 1 s007
rlabel pdcontact 2535 1 2537 2 1 s010
rlabel ndcontact 2535 -42 2537 -41 1 s011
rlabel metal1 2512 -22 2515 -21 1 s0_q
rlabel metal1 2475 -22 2479 -21 1 s009
rlabel metal1 2366 -22 2369 -21 1 s004
rlabel metal1 2329 -22 2333 -21 1 s003
rlabel pdcontact 2013 102 2015 103 1 s301
rlabel ndcontact 2013 59 2015 60 1 s302
rlabel pdcontact 2091 102 2093 103 1 s305
rlabel ndcontact 2091 59 2093 60 1 s306
rlabel ndcontact 2159 59 2161 60 1 s308
rlabel pdcontact 2159 102 2161 103 1 s307
rlabel pdcontact 2237 102 2239 103 1 s310
rlabel ndcontact 2237 59 2239 60 1 s311
rlabel metal1 2214 79 2217 80 1 s3_q
rlabel metal1 2177 79 2181 80 1 s309
rlabel metal1 2068 79 2071 80 1 s304
rlabel metal1 2031 79 2035 80 1 s303
rlabel metal1 1996 79 1999 80 1 s3
rlabel metal1 1995 86 1997 87 1 clks3
rlabel metal1 1995 72 1997 73 1 clks3_bar
rlabel metal1 2294 79 2297 80 1 s1
rlabel metal1 2293 72 2295 73 1 clks1_bar
rlabel metal1 2293 86 2295 87 1 clks1
rlabel ndcontact 2311 59 2313 60 1 s102
rlabel pdcontact 2311 102 2313 103 1 s101
rlabel pdcontact 2389 102 2391 103 1 s105
rlabel ndcontact 2389 59 2391 60 1 s106
rlabel pdcontact 2457 102 2459 103 1 s107
rlabel ndcontact 2457 59 2459 60 1 s108
rlabel pdcontact 2535 102 2537 103 1 s110
rlabel ndcontact 2535 59 2537 60 1 s111
rlabel metal1 2512 79 2515 80 1 s1_q
rlabel metal1 2475 79 2479 80 1 s109
rlabel metal1 2366 79 2369 80 1 s104
rlabel metal1 2329 79 2333 80 1 s103
rlabel metal1 2043 161 2047 162 1 gnd
rlabel metal1 2039 198 2050 199 5 vdd
rlabel metal1 2189 161 2193 162 1 gnd
rlabel metal1 2185 198 2196 199 5 vdd
rlabel metal1 1988 169 1990 170 1 clkc4_bar
rlabel metal1 1988 183 1990 184 1 clkc4
rlabel metal1 1989 176 1992 177 1 c4
rlabel ndcontact 2006 156 2008 157 1 c402
rlabel pdcontact 2006 199 2008 200 1 c401
rlabel metal1 2024 176 2028 177 1 c403
rlabel metal1 2061 176 2064 177 1 c404
rlabel pdcontact 2084 199 2086 200 1 c405
rlabel ndcontact 2084 156 2086 157 1 c406
rlabel ndcontact 2152 156 2154 157 1 c408
rlabel pdcontact 2152 199 2154 200 1 c407
rlabel metal1 2170 176 2174 177 1 c409
rlabel metal1 2207 176 2210 177 1 c4_q
rlabel pdcontact 2230 199 2232 200 1 c410
rlabel ndcontact 2230 156 2232 157 1 c411
rlabel metal1 911 -37 915 -36 1 gnd
rlabel metal1 907 0 918 1 5 vdd
rlabel metal1 759 -37 763 -36 1 gnd
rlabel metal1 755 0 766 1 5 vdd
rlabel metal1 613 -37 617 -36 1 gnd
rlabel metal1 609 0 620 1 5 vdd
rlabel metal1 461 -37 465 -36 1 gnd
rlabel metal1 457 0 468 1 5 vdd
rlabel metal1 315 -37 319 -36 1 gnd
rlabel metal1 311 0 322 1 5 vdd
rlabel metal1 163 -37 167 -36 1 gnd
rlabel metal1 159 0 170 1 5 vdd
<< end >>

magic
tech scmos
timestamp 1619385914
<< nwell >>
rect -65 -2 -33 18
rect -6 -28 26 14
rect -76 -59 -22 -39
<< ntransistor >>
rect -58 -21 -56 -17
rect -42 -21 -40 -17
rect 5 -46 7 -42
rect 13 -46 15 -42
rect -65 -69 -63 -65
rect -35 -69 -33 -65
rect 5 -68 7 -64
rect 13 -68 15 -64
<< ptransistor >>
rect -54 4 -52 12
rect -46 4 -44 12
rect 5 0 7 8
rect 13 0 15 8
rect 5 -22 7 -14
rect 13 -22 15 -14
rect -65 -53 -63 -45
rect -35 -53 -33 -45
<< ndiffusion >>
rect -59 -21 -58 -17
rect -56 -21 -55 -17
rect -43 -21 -42 -17
rect -40 -21 -39 -17
rect 4 -46 5 -42
rect 7 -46 8 -42
rect 12 -46 13 -42
rect 15 -46 16 -42
rect -66 -69 -65 -65
rect -63 -69 -62 -65
rect -36 -69 -35 -65
rect -33 -69 -32 -65
rect 4 -68 5 -64
rect 7 -68 8 -64
rect 12 -68 13 -64
rect 15 -68 16 -64
<< pdiffusion >>
rect -55 4 -54 12
rect -52 4 -51 12
rect -47 4 -46 12
rect -44 4 -43 12
rect 4 0 5 8
rect 7 0 8 8
rect 12 0 13 8
rect 15 0 16 8
rect 4 -22 5 -14
rect 7 -22 8 -14
rect 12 -22 13 -14
rect 15 -22 16 -14
rect -66 -53 -65 -45
rect -63 -53 -62 -45
rect -36 -53 -35 -45
rect -33 -53 -32 -45
<< ndcontact >>
rect -63 -21 -59 -17
rect -55 -21 -51 -17
rect -47 -21 -43 -17
rect -39 -21 -35 -17
rect 0 -46 4 -42
rect 8 -46 12 -42
rect 16 -46 20 -42
rect -70 -69 -66 -65
rect -62 -69 -58 -65
rect -40 -69 -36 -65
rect -32 -69 -28 -65
rect 0 -68 4 -64
rect 8 -68 12 -64
rect 16 -68 20 -64
<< pdcontact >>
rect -59 4 -55 12
rect -51 4 -47 12
rect -43 4 -39 12
rect 0 0 4 8
rect 8 0 12 8
rect 16 0 20 8
rect 0 -22 4 -14
rect 8 -22 12 -14
rect 16 -22 20 -14
rect -70 -53 -66 -45
rect -62 -53 -58 -45
rect -40 -53 -36 -45
rect -32 -53 -28 -45
<< polysilicon >>
rect -54 12 -52 15
rect -46 12 -44 15
rect 5 8 7 11
rect 13 8 15 11
rect -54 3 -52 4
rect -58 1 -52 3
rect -46 3 -44 4
rect -46 1 -40 3
rect -58 -17 -56 1
rect -42 -17 -40 1
rect 5 -7 7 0
rect 13 -7 15 0
rect 5 -14 7 -11
rect 13 -14 15 -11
rect -58 -24 -56 -21
rect -42 -24 -40 -21
rect 5 -42 7 -22
rect 13 -30 15 -22
rect 13 -42 15 -34
rect -65 -45 -63 -42
rect -35 -45 -33 -42
rect 5 -49 7 -46
rect 13 -49 15 -46
rect -65 -65 -63 -53
rect -35 -65 -33 -53
rect 5 -64 7 -57
rect 13 -64 15 -57
rect -65 -72 -63 -69
rect -35 -72 -33 -69
rect 5 -71 7 -68
rect 13 -71 15 -68
<< polycontact >>
rect -62 -3 -58 1
rect -46 -7 -42 -3
rect 1 -7 5 -3
rect 15 -7 19 -3
rect 1 -36 5 -32
rect 15 -29 19 -25
rect 15 -39 19 -35
rect -69 -61 -65 -57
rect -39 -61 -35 -57
rect 1 -61 5 -57
rect 15 -61 19 -57
<< metal1 >>
rect -87 24 56 27
rect -75 -38 -71 24
rect -59 12 -55 24
rect -63 -3 -62 1
rect -47 -7 -46 -3
rect -39 -11 -35 12
rect -55 -14 -35 -11
rect -55 -17 -51 -14
rect -39 -17 -35 -14
rect -18 -14 -14 24
rect 0 8 4 24
rect 20 2 43 6
rect -2 -7 1 -3
rect 19 -7 22 -3
rect -18 -18 0 -14
rect -63 -25 -59 -21
rect -47 -25 -43 -21
rect 39 -16 43 2
rect 20 -20 43 -16
rect 47 -15 51 15
rect 47 -19 56 -15
rect -63 -28 -14 -25
rect -75 -41 -36 -38
rect -87 -48 -82 -44
rect -70 -45 -66 -41
rect -40 -45 -36 -41
rect -18 -42 -14 -28
rect 19 -29 22 -25
rect 39 -30 43 -20
rect -3 -36 1 -32
rect 39 -34 56 -30
rect 19 -39 22 -35
rect 39 -42 43 -34
rect -62 -56 -58 -53
rect -87 -61 -78 -57
rect -73 -61 -69 -57
rect -62 -65 -58 -61
rect -42 -61 -39 -57
rect -32 -65 -28 -53
rect -18 -46 0 -42
rect 20 -46 43 -42
rect -70 -83 -66 -69
rect -40 -83 -36 -69
rect -18 -83 -14 -46
rect 1 -57 5 -55
rect 15 -57 19 -55
rect 39 -64 43 -46
rect 20 -68 43 -64
rect 0 -83 4 -68
rect -87 -86 56 -83
<< m2contact >>
rect -52 -8 -47 -3
rect 22 -30 27 -25
rect -8 -36 -3 -31
rect -78 -62 -73 -57
rect -28 -62 -23 -57
rect 15 -55 20 -50
<< metal2 >>
rect -23 14 38 18
rect -51 -29 -47 -8
rect -23 -29 -19 14
rect 34 -25 38 14
rect -51 -32 -19 -29
rect 27 -29 38 -25
rect -23 -62 -19 -32
rect -77 -73 -73 -62
rect -8 -73 -4 -36
rect 34 -51 38 -29
rect 20 -55 38 -51
rect -77 -77 -4 -73
<< m123contact >>
rect -68 -4 -63 1
rect -35 -13 -30 -8
rect -7 -8 -2 -3
rect 22 -8 27 -3
rect 42 10 47 15
rect -82 -49 -77 -44
rect -62 -61 -57 -56
rect -47 -62 -42 -57
rect 22 -39 27 -34
rect 0 -55 5 -50
<< metal3 >>
rect -30 19 47 23
rect -68 -33 -64 -4
rect -30 -13 -26 19
rect 42 15 47 19
rect -13 -8 -7 -3
rect 27 -8 33 -4
rect -13 -33 -9 -8
rect -68 -37 -9 -33
rect 29 -34 33 -8
rect -82 -78 -79 -49
rect -55 -56 -51 -37
rect -13 -50 -9 -37
rect 27 -39 33 -34
rect -13 -55 0 -50
rect -57 -60 -51 -56
rect -47 -78 -43 -62
rect 23 -78 27 -39
rect -82 -82 27 -78
<< labels >>
rlabel metal1 -86 -60 -84 -59 3 a0
rlabel metal1 -86 -47 -84 -46 3 b0
rlabel metal1 -60 -64 -59 -63 1 a0_bar
rlabel metal1 -30 -64 -29 -63 1 b0_bar
rlabel pdcontact -49 6 -48 7 1 an0
rlabel pdcontact 9 3 10 4 1 xr00
rlabel pdcontact 9 -19 10 -18 1 xr01
rlabel ndcontact 9 -45 10 -44 1 xr02
rlabel ndcontact 9 -67 10 -66 1 xr03
rlabel metal1 50 -18 52 -17 1 g0
rlabel metal1 50 -33 52 -32 1 p0
rlabel metal1 -17 -85 -15 -84 1 gnd
rlabel metal1 -17 25 -15 26 5 vdd
<< end >>

magic
tech scmos
timestamp 1619418083
<< nwell >>
rect -47 -2 -15 18
rect 12 -28 44 14
rect 124 -2 156 18
rect 183 -28 215 14
rect -58 -59 -4 -39
rect 113 -59 167 -39
rect -47 -121 -15 -101
rect 12 -147 44 -105
rect 124 -121 156 -101
rect 183 -147 215 -105
rect -58 -178 -4 -158
rect 113 -178 167 -158
<< ntransistor >>
rect -40 -21 -38 -17
rect -24 -21 -22 -17
rect 131 -21 133 -17
rect 147 -21 149 -17
rect 23 -46 25 -42
rect 31 -46 33 -42
rect 194 -46 196 -42
rect 202 -46 204 -42
rect -47 -69 -45 -65
rect -17 -69 -15 -65
rect 23 -68 25 -64
rect 31 -68 33 -64
rect 124 -69 126 -65
rect 154 -69 156 -65
rect 194 -68 196 -64
rect 202 -68 204 -64
rect -40 -140 -38 -136
rect -24 -140 -22 -136
rect 131 -140 133 -136
rect 147 -140 149 -136
rect 23 -165 25 -161
rect 31 -165 33 -161
rect 194 -165 196 -161
rect 202 -165 204 -161
rect -47 -188 -45 -184
rect -17 -188 -15 -184
rect 23 -187 25 -183
rect 31 -187 33 -183
rect 124 -188 126 -184
rect 154 -188 156 -184
rect 194 -187 196 -183
rect 202 -187 204 -183
<< ptransistor >>
rect -36 4 -34 12
rect -28 4 -26 12
rect 23 0 25 8
rect 31 0 33 8
rect 135 4 137 12
rect 143 4 145 12
rect 23 -22 25 -14
rect 31 -22 33 -14
rect 194 0 196 8
rect 202 0 204 8
rect 194 -22 196 -14
rect 202 -22 204 -14
rect -47 -53 -45 -45
rect -17 -53 -15 -45
rect 124 -53 126 -45
rect 154 -53 156 -45
rect -36 -115 -34 -107
rect -28 -115 -26 -107
rect 23 -119 25 -111
rect 31 -119 33 -111
rect 135 -115 137 -107
rect 143 -115 145 -107
rect 23 -141 25 -133
rect 31 -141 33 -133
rect 194 -119 196 -111
rect 202 -119 204 -111
rect 194 -141 196 -133
rect 202 -141 204 -133
rect -47 -172 -45 -164
rect -17 -172 -15 -164
rect 124 -172 126 -164
rect 154 -172 156 -164
<< ndiffusion >>
rect -41 -21 -40 -17
rect -38 -21 -37 -17
rect -25 -21 -24 -17
rect -22 -21 -21 -17
rect 130 -21 131 -17
rect 133 -21 134 -17
rect 146 -21 147 -17
rect 149 -21 150 -17
rect 22 -46 23 -42
rect 25 -46 26 -42
rect 30 -46 31 -42
rect 33 -46 34 -42
rect 193 -46 194 -42
rect 196 -46 197 -42
rect 201 -46 202 -42
rect 204 -46 205 -42
rect -48 -69 -47 -65
rect -45 -69 -44 -65
rect -18 -69 -17 -65
rect -15 -69 -14 -65
rect 22 -68 23 -64
rect 25 -68 26 -64
rect 30 -68 31 -64
rect 33 -68 34 -64
rect 123 -69 124 -65
rect 126 -69 127 -65
rect 153 -69 154 -65
rect 156 -69 157 -65
rect 193 -68 194 -64
rect 196 -68 197 -64
rect 201 -68 202 -64
rect 204 -68 205 -64
rect -41 -140 -40 -136
rect -38 -140 -37 -136
rect -25 -140 -24 -136
rect -22 -140 -21 -136
rect 130 -140 131 -136
rect 133 -140 134 -136
rect 146 -140 147 -136
rect 149 -140 150 -136
rect 22 -165 23 -161
rect 25 -165 26 -161
rect 30 -165 31 -161
rect 33 -165 34 -161
rect 193 -165 194 -161
rect 196 -165 197 -161
rect 201 -165 202 -161
rect 204 -165 205 -161
rect -48 -188 -47 -184
rect -45 -188 -44 -184
rect -18 -188 -17 -184
rect -15 -188 -14 -184
rect 22 -187 23 -183
rect 25 -187 26 -183
rect 30 -187 31 -183
rect 33 -187 34 -183
rect 123 -188 124 -184
rect 126 -188 127 -184
rect 153 -188 154 -184
rect 156 -188 157 -184
rect 193 -187 194 -183
rect 196 -187 197 -183
rect 201 -187 202 -183
rect 204 -187 205 -183
<< pdiffusion >>
rect -37 4 -36 12
rect -34 4 -33 12
rect -29 4 -28 12
rect -26 4 -25 12
rect 22 0 23 8
rect 25 0 26 8
rect 30 0 31 8
rect 33 0 34 8
rect 134 4 135 12
rect 137 4 138 12
rect 142 4 143 12
rect 145 4 146 12
rect 22 -22 23 -14
rect 25 -22 26 -14
rect 30 -22 31 -14
rect 33 -22 34 -14
rect 193 0 194 8
rect 196 0 197 8
rect 201 0 202 8
rect 204 0 205 8
rect 193 -22 194 -14
rect 196 -22 197 -14
rect 201 -22 202 -14
rect 204 -22 205 -14
rect -48 -53 -47 -45
rect -45 -53 -44 -45
rect -18 -53 -17 -45
rect -15 -53 -14 -45
rect 123 -53 124 -45
rect 126 -53 127 -45
rect 153 -53 154 -45
rect 156 -53 157 -45
rect -37 -115 -36 -107
rect -34 -115 -33 -107
rect -29 -115 -28 -107
rect -26 -115 -25 -107
rect 22 -119 23 -111
rect 25 -119 26 -111
rect 30 -119 31 -111
rect 33 -119 34 -111
rect 134 -115 135 -107
rect 137 -115 138 -107
rect 142 -115 143 -107
rect 145 -115 146 -107
rect 22 -141 23 -133
rect 25 -141 26 -133
rect 30 -141 31 -133
rect 33 -141 34 -133
rect 193 -119 194 -111
rect 196 -119 197 -111
rect 201 -119 202 -111
rect 204 -119 205 -111
rect 193 -141 194 -133
rect 196 -141 197 -133
rect 201 -141 202 -133
rect 204 -141 205 -133
rect -48 -172 -47 -164
rect -45 -172 -44 -164
rect -18 -172 -17 -164
rect -15 -172 -14 -164
rect 123 -172 124 -164
rect 126 -172 127 -164
rect 153 -172 154 -164
rect 156 -172 157 -164
<< ndcontact >>
rect -45 -21 -41 -17
rect -37 -21 -33 -17
rect -29 -21 -25 -17
rect -21 -21 -17 -17
rect 126 -21 130 -17
rect 134 -21 138 -17
rect 142 -21 146 -17
rect 150 -21 154 -17
rect 18 -46 22 -42
rect 26 -46 30 -42
rect 34 -46 38 -42
rect 189 -46 193 -42
rect 197 -46 201 -42
rect 205 -46 209 -42
rect -52 -69 -48 -65
rect -44 -69 -40 -65
rect -22 -69 -18 -65
rect -14 -69 -10 -65
rect 18 -68 22 -64
rect 26 -68 30 -64
rect 34 -68 38 -64
rect 119 -69 123 -65
rect 127 -69 131 -65
rect 149 -69 153 -65
rect 157 -69 161 -65
rect 189 -68 193 -64
rect 197 -68 201 -64
rect 205 -68 209 -64
rect -45 -140 -41 -136
rect -37 -140 -33 -136
rect -29 -140 -25 -136
rect -21 -140 -17 -136
rect 126 -140 130 -136
rect 134 -140 138 -136
rect 142 -140 146 -136
rect 150 -140 154 -136
rect 18 -165 22 -161
rect 26 -165 30 -161
rect 34 -165 38 -161
rect 189 -165 193 -161
rect 197 -165 201 -161
rect 205 -165 209 -161
rect -52 -188 -48 -184
rect -44 -188 -40 -184
rect -22 -188 -18 -184
rect -14 -188 -10 -184
rect 18 -187 22 -183
rect 26 -187 30 -183
rect 34 -187 38 -183
rect 119 -188 123 -184
rect 127 -188 131 -184
rect 149 -188 153 -184
rect 157 -188 161 -184
rect 189 -187 193 -183
rect 197 -187 201 -183
rect 205 -187 209 -183
<< pdcontact >>
rect -41 4 -37 12
rect -33 4 -29 12
rect -25 4 -21 12
rect 18 0 22 8
rect 26 0 30 8
rect 34 0 38 8
rect 130 4 134 12
rect 138 4 142 12
rect 146 4 150 12
rect 18 -22 22 -14
rect 26 -22 30 -14
rect 34 -22 38 -14
rect 189 0 193 8
rect 197 0 201 8
rect 205 0 209 8
rect 189 -22 193 -14
rect 197 -22 201 -14
rect 205 -22 209 -14
rect -52 -53 -48 -45
rect -44 -53 -40 -45
rect -22 -53 -18 -45
rect -14 -53 -10 -45
rect 119 -53 123 -45
rect 127 -53 131 -45
rect 149 -53 153 -45
rect 157 -53 161 -45
rect -41 -115 -37 -107
rect -33 -115 -29 -107
rect -25 -115 -21 -107
rect 18 -119 22 -111
rect 26 -119 30 -111
rect 34 -119 38 -111
rect 130 -115 134 -107
rect 138 -115 142 -107
rect 146 -115 150 -107
rect 18 -141 22 -133
rect 26 -141 30 -133
rect 34 -141 38 -133
rect 189 -119 193 -111
rect 197 -119 201 -111
rect 205 -119 209 -111
rect 189 -141 193 -133
rect 197 -141 201 -133
rect 205 -141 209 -133
rect -52 -172 -48 -164
rect -44 -172 -40 -164
rect -22 -172 -18 -164
rect -14 -172 -10 -164
rect 119 -172 123 -164
rect 127 -172 131 -164
rect 149 -172 153 -164
rect 157 -172 161 -164
<< polysilicon >>
rect -36 12 -34 15
rect -28 12 -26 15
rect 135 12 137 15
rect 143 12 145 15
rect 23 8 25 11
rect 31 8 33 11
rect -36 3 -34 4
rect -40 1 -34 3
rect -28 3 -26 4
rect -28 1 -22 3
rect -40 -17 -38 1
rect -24 -17 -22 1
rect 194 8 196 11
rect 202 8 204 11
rect 135 3 137 4
rect 131 1 137 3
rect 143 3 145 4
rect 143 1 149 3
rect 23 -7 25 0
rect 31 -7 33 0
rect 23 -14 25 -11
rect 31 -14 33 -11
rect -40 -24 -38 -21
rect -24 -24 -22 -21
rect 131 -17 133 1
rect 147 -17 149 1
rect 194 -7 196 0
rect 202 -7 204 0
rect 194 -14 196 -11
rect 202 -14 204 -11
rect 23 -42 25 -22
rect 31 -30 33 -22
rect 131 -24 133 -21
rect 147 -24 149 -21
rect 31 -42 33 -34
rect 194 -42 196 -22
rect 202 -30 204 -22
rect 202 -42 204 -34
rect -47 -45 -45 -42
rect -17 -45 -15 -42
rect 124 -45 126 -42
rect 154 -45 156 -42
rect 23 -49 25 -46
rect 31 -49 33 -46
rect 194 -49 196 -46
rect 202 -49 204 -46
rect -47 -65 -45 -53
rect -17 -65 -15 -53
rect 23 -64 25 -57
rect 31 -64 33 -57
rect 124 -65 126 -53
rect 154 -65 156 -53
rect 194 -64 196 -57
rect 202 -64 204 -57
rect -47 -72 -45 -69
rect -17 -72 -15 -69
rect 23 -71 25 -68
rect 31 -71 33 -68
rect 124 -72 126 -69
rect 154 -72 156 -69
rect 194 -71 196 -68
rect 202 -71 204 -68
rect -36 -107 -34 -104
rect -28 -107 -26 -104
rect 135 -107 137 -104
rect 143 -107 145 -104
rect 23 -111 25 -108
rect 31 -111 33 -108
rect -36 -116 -34 -115
rect -40 -118 -34 -116
rect -28 -116 -26 -115
rect -28 -118 -22 -116
rect -40 -136 -38 -118
rect -24 -136 -22 -118
rect 194 -111 196 -108
rect 202 -111 204 -108
rect 135 -116 137 -115
rect 131 -118 137 -116
rect 143 -116 145 -115
rect 143 -118 149 -116
rect 23 -126 25 -119
rect 31 -126 33 -119
rect 23 -133 25 -130
rect 31 -133 33 -130
rect -40 -143 -38 -140
rect -24 -143 -22 -140
rect 131 -136 133 -118
rect 147 -136 149 -118
rect 194 -126 196 -119
rect 202 -126 204 -119
rect 194 -133 196 -130
rect 202 -133 204 -130
rect 23 -161 25 -141
rect 31 -149 33 -141
rect 131 -143 133 -140
rect 147 -143 149 -140
rect 31 -161 33 -153
rect 194 -161 196 -141
rect 202 -149 204 -141
rect 202 -161 204 -153
rect -47 -164 -45 -161
rect -17 -164 -15 -161
rect 124 -164 126 -161
rect 154 -164 156 -161
rect 23 -168 25 -165
rect 31 -168 33 -165
rect 194 -168 196 -165
rect 202 -168 204 -165
rect -47 -184 -45 -172
rect -17 -184 -15 -172
rect 23 -183 25 -176
rect 31 -183 33 -176
rect 124 -184 126 -172
rect 154 -184 156 -172
rect 194 -183 196 -176
rect 202 -183 204 -176
rect -47 -191 -45 -188
rect -17 -191 -15 -188
rect 23 -190 25 -187
rect 31 -190 33 -187
rect 124 -191 126 -188
rect 154 -191 156 -188
rect 194 -190 196 -187
rect 202 -190 204 -187
<< polycontact >>
rect -44 -3 -40 1
rect -28 -7 -24 -3
rect 19 -7 23 -3
rect 127 -3 131 1
rect 33 -7 37 -3
rect 143 -7 147 -3
rect 190 -7 194 -3
rect 204 -7 208 -3
rect 19 -36 23 -32
rect 33 -29 37 -25
rect 33 -39 37 -35
rect 190 -36 194 -32
rect 204 -29 208 -25
rect 204 -39 208 -35
rect -51 -61 -47 -57
rect -21 -61 -17 -57
rect 19 -61 23 -57
rect 33 -61 37 -57
rect 120 -61 124 -57
rect 150 -61 154 -57
rect 190 -61 194 -57
rect 204 -61 208 -57
rect -44 -122 -40 -118
rect -28 -126 -24 -122
rect 19 -126 23 -122
rect 127 -122 131 -118
rect 33 -126 37 -122
rect 143 -126 147 -122
rect 190 -126 194 -122
rect 204 -126 208 -122
rect 19 -155 23 -151
rect 33 -148 37 -144
rect 33 -158 37 -154
rect 190 -155 194 -151
rect 204 -148 208 -144
rect 204 -158 208 -154
rect -51 -180 -47 -176
rect -21 -180 -17 -176
rect 19 -180 23 -176
rect 33 -180 37 -176
rect 120 -180 124 -176
rect 150 -180 154 -176
rect 190 -180 194 -176
rect 204 -180 208 -176
<< metal1 >>
rect -91 59 -45 63
rect -91 50 -52 54
rect -91 41 -64 45
rect -91 32 -82 36
rect -56 36 -52 50
rect -49 45 -45 59
rect 245 58 265 62
rect 254 49 265 53
rect -49 41 107 45
rect 131 41 265 45
rect -56 32 89 36
rect 122 32 265 36
rect -91 24 265 27
rect -77 -92 -73 24
rect -57 -38 -53 24
rect -41 12 -37 24
rect -45 -3 -44 1
rect -29 -7 -28 -3
rect -21 -11 -17 12
rect -37 -14 -17 -11
rect -37 -17 -33 -14
rect -21 -17 -17 -14
rect 0 -14 4 24
rect 18 8 22 24
rect 38 2 61 6
rect 16 -7 19 -3
rect 37 -7 40 -3
rect 0 -18 18 -14
rect -45 -25 -41 -21
rect -29 -25 -25 -21
rect 57 -16 61 2
rect 38 -20 61 -16
rect -45 -28 4 -25
rect -57 -41 -18 -38
rect -69 -48 -64 -44
rect -52 -45 -48 -41
rect -22 -45 -18 -41
rect 0 -42 4 -28
rect 37 -29 40 -25
rect 57 -30 61 -20
rect 15 -36 19 -32
rect 57 -34 70 -30
rect 37 -39 40 -35
rect 57 -42 61 -34
rect -44 -56 -40 -53
rect -69 -61 -60 -57
rect -55 -61 -51 -57
rect -44 -65 -40 -61
rect -24 -61 -21 -57
rect -14 -65 -10 -53
rect 0 -46 18 -42
rect 38 -46 61 -42
rect -52 -83 -48 -69
rect -22 -83 -18 -69
rect 0 -83 4 -46
rect 19 -57 23 -55
rect 33 -57 37 -55
rect 57 -64 61 -46
rect 38 -68 61 -64
rect 18 -83 22 -68
rect -64 -86 22 -83
rect -77 -95 22 -92
rect -57 -157 -53 -95
rect -41 -107 -37 -95
rect -45 -122 -44 -118
rect -29 -126 -28 -122
rect -21 -130 -17 -107
rect -37 -133 -17 -130
rect -37 -136 -33 -133
rect -21 -136 -17 -133
rect 0 -133 4 -95
rect 18 -111 22 -95
rect 64 -104 68 -92
rect 38 -117 61 -113
rect 16 -126 19 -122
rect 37 -126 40 -122
rect 0 -137 18 -133
rect -45 -144 -41 -140
rect -29 -144 -25 -140
rect 57 -135 61 -117
rect 38 -139 61 -135
rect -45 -147 4 -144
rect -57 -160 -18 -157
rect -69 -167 -64 -163
rect -52 -164 -48 -160
rect -22 -164 -18 -160
rect 0 -161 4 -147
rect 37 -148 40 -144
rect 57 -149 61 -139
rect 79 -149 83 15
rect 94 -92 98 24
rect 114 -38 118 24
rect 130 12 134 24
rect 126 -3 127 1
rect 142 -7 143 -3
rect 150 -11 154 12
rect 134 -14 154 -11
rect 134 -17 138 -14
rect 150 -17 154 -14
rect 171 -14 175 24
rect 189 8 193 24
rect 209 2 232 6
rect 187 -7 190 -3
rect 208 -7 211 -3
rect 171 -18 189 -14
rect 126 -25 130 -21
rect 142 -25 146 -21
rect 228 -16 232 2
rect 209 -20 232 -16
rect 126 -28 175 -25
rect 114 -41 153 -38
rect 102 -48 107 -44
rect 119 -45 123 -41
rect 149 -45 153 -41
rect 171 -42 175 -28
rect 208 -29 211 -25
rect 228 -30 232 -20
rect 240 -30 244 13
rect 186 -36 190 -32
rect 228 -34 244 -30
rect 208 -39 211 -35
rect 228 -42 232 -34
rect 127 -56 131 -53
rect 102 -61 111 -57
rect 116 -61 120 -57
rect 127 -65 131 -61
rect 147 -61 150 -57
rect 157 -65 161 -53
rect 171 -46 189 -42
rect 209 -46 232 -42
rect 119 -83 123 -69
rect 149 -83 153 -69
rect 171 -83 175 -46
rect 190 -57 194 -55
rect 204 -57 208 -55
rect 228 -64 232 -46
rect 209 -68 232 -64
rect 189 -83 193 -68
rect 107 -86 193 -83
rect 94 -95 193 -92
rect 15 -155 19 -151
rect 57 -153 83 -149
rect 37 -158 40 -154
rect 57 -161 61 -153
rect 114 -157 118 -95
rect 130 -107 134 -95
rect 126 -122 127 -118
rect 142 -126 143 -122
rect 150 -130 154 -107
rect 134 -133 154 -130
rect 134 -136 138 -133
rect 150 -136 154 -133
rect 171 -133 175 -95
rect 189 -111 193 -95
rect 234 -104 238 -92
rect 209 -117 232 -113
rect 187 -126 190 -122
rect 208 -126 211 -122
rect 171 -137 189 -133
rect 126 -144 130 -140
rect 142 -144 146 -140
rect 228 -135 232 -117
rect 209 -139 232 -135
rect 126 -147 175 -144
rect 114 -160 153 -157
rect -44 -175 -40 -172
rect -69 -180 -60 -176
rect -55 -180 -51 -176
rect -44 -184 -40 -180
rect -24 -180 -21 -176
rect -14 -184 -10 -172
rect 0 -165 18 -161
rect 38 -165 61 -161
rect -91 -205 -74 -202
rect -52 -202 -48 -188
rect -22 -202 -18 -188
rect 0 -202 4 -165
rect 19 -176 23 -174
rect 33 -176 37 -174
rect 57 -183 61 -165
rect 102 -167 107 -163
rect 119 -164 123 -160
rect 149 -164 153 -160
rect 171 -161 175 -147
rect 208 -148 211 -144
rect 228 -149 232 -139
rect 250 -149 254 13
rect 186 -155 190 -151
rect 228 -153 254 -149
rect 208 -158 211 -154
rect 228 -161 232 -153
rect 127 -175 131 -172
rect 102 -180 111 -176
rect 116 -180 120 -176
rect 38 -187 61 -183
rect 127 -184 131 -180
rect 147 -180 150 -176
rect 157 -184 161 -172
rect 171 -165 189 -161
rect 209 -165 232 -161
rect 18 -202 22 -187
rect -69 -205 97 -202
rect 119 -202 123 -188
rect 149 -202 153 -188
rect 171 -202 175 -165
rect 190 -176 194 -174
rect 204 -176 208 -174
rect 228 -183 232 -165
rect 209 -187 232 -183
rect 189 -202 193 -187
rect 102 -205 266 -202
rect -91 -214 -59 -210
rect -51 -214 112 -210
rect 120 -214 266 -210
rect -91 -223 -85 -219
rect -51 -228 -46 -214
rect -91 -232 -46 -228
rect -42 -223 84 -219
rect -42 -237 -38 -223
rect 120 -228 124 -214
rect 78 -232 124 -228
rect 128 -223 266 -219
rect -91 -241 -38 -237
rect 128 -237 132 -223
rect 248 -232 266 -228
rect 69 -241 132 -237
rect 239 -241 266 -237
<< m2contact >>
rect 240 57 245 62
rect 249 49 254 54
rect 126 41 131 46
rect 117 32 122 37
rect -34 -8 -29 -3
rect 79 15 84 20
rect 40 -30 45 -25
rect 10 -36 15 -31
rect 70 -34 75 -29
rect -60 -62 -55 -57
rect -10 -62 -5 -57
rect 33 -55 38 -50
rect -69 -88 -64 -83
rect -34 -127 -29 -122
rect 40 -149 45 -144
rect 137 -8 142 -3
rect 240 13 245 18
rect 249 13 254 18
rect 211 -30 216 -25
rect 181 -36 186 -31
rect 111 -62 116 -57
rect 161 -62 166 -57
rect 204 -55 209 -50
rect 102 -88 107 -83
rect 10 -155 15 -150
rect 137 -127 142 -122
rect -60 -181 -55 -176
rect -10 -181 -5 -176
rect -74 -205 -69 -200
rect 33 -174 38 -169
rect 211 -149 216 -144
rect 181 -155 186 -150
rect 111 -181 116 -176
rect 161 -181 166 -176
rect 97 -205 102 -200
rect 204 -174 209 -169
rect -59 -214 -54 -209
rect 112 -214 117 -209
rect -85 -223 -80 -218
rect 84 -223 89 -218
<< metal2 >>
rect 71 58 130 62
rect -5 14 56 18
rect -33 -29 -29 -8
rect -5 -29 -1 14
rect 52 -25 56 14
rect -33 -32 -1 -29
rect 45 -29 56 -25
rect 71 -29 75 58
rect 79 50 121 54
rect 79 20 83 50
rect 117 37 121 50
rect 126 46 130 58
rect 240 18 244 57
rect 250 18 254 49
rect 166 14 227 18
rect -5 -62 -1 -32
rect -59 -73 -55 -62
rect 10 -73 14 -36
rect 52 -51 56 -29
rect 138 -29 142 -8
rect 166 -29 170 14
rect 223 -25 227 14
rect 138 -32 170 -29
rect 216 -29 227 -25
rect 38 -55 56 -51
rect 166 -62 170 -32
rect 112 -73 116 -62
rect 181 -73 185 -36
rect 223 -51 227 -29
rect 209 -55 227 -51
rect -87 -77 14 -73
rect 84 -77 185 -73
rect -87 -111 -83 -77
rect -69 -97 -65 -88
rect -77 -101 -65 -97
rect -87 -114 -81 -111
rect -85 -218 -81 -114
rect -77 -197 -73 -101
rect -5 -105 56 -101
rect -33 -148 -29 -127
rect -5 -148 -1 -105
rect 52 -144 56 -105
rect -33 -151 -1 -148
rect 45 -148 56 -144
rect -5 -181 -1 -151
rect -59 -192 -55 -181
rect 10 -192 14 -155
rect 52 -170 56 -148
rect 38 -174 56 -170
rect -59 -196 14 -192
rect -77 -200 -69 -197
rect -59 -209 -55 -196
rect 84 -218 88 -77
rect 102 -97 106 -88
rect 94 -101 106 -97
rect 94 -197 98 -101
rect 166 -105 227 -101
rect 138 -148 142 -127
rect 166 -148 170 -105
rect 223 -144 227 -105
rect 138 -151 170 -148
rect 216 -148 227 -144
rect 166 -181 170 -151
rect 112 -192 116 -181
rect 181 -192 185 -155
rect 223 -170 227 -148
rect 209 -174 227 -170
rect 112 -196 185 -192
rect 94 -200 102 -197
rect 112 -209 116 -196
<< m123contact >>
rect -64 41 -59 46
rect -82 32 -77 37
rect -50 -4 -45 1
rect -17 -13 -12 -8
rect 11 -8 16 -3
rect 40 -8 45 -3
rect 107 41 112 46
rect 89 32 94 37
rect 121 -4 126 1
rect -64 -49 -59 -44
rect -44 -61 -39 -56
rect -29 -62 -24 -57
rect 40 -39 45 -34
rect 18 -55 23 -50
rect 154 -13 159 -8
rect 182 -8 187 -3
rect 211 -8 216 -3
rect 107 -49 112 -44
rect 127 -61 132 -56
rect 142 -62 147 -57
rect 211 -39 216 -34
rect 189 -55 194 -50
rect 64 -92 69 -87
rect -50 -123 -45 -118
rect -17 -132 -12 -127
rect 11 -127 16 -122
rect 40 -127 45 -122
rect 64 -109 69 -104
rect -64 -168 -59 -163
rect -44 -180 -39 -175
rect -29 -181 -24 -176
rect 40 -158 45 -153
rect 18 -174 23 -169
rect 234 -92 239 -87
rect 121 -123 126 -118
rect 154 -132 159 -127
rect 182 -127 187 -122
rect 211 -127 216 -122
rect 234 -109 239 -104
rect 107 -168 112 -163
rect 127 -180 132 -175
rect 142 -181 147 -176
rect 211 -158 216 -153
rect 189 -174 194 -169
rect 73 -232 78 -227
rect 243 -233 248 -228
rect 64 -241 69 -236
rect 234 -241 239 -236
<< metal3 >>
rect -82 -105 -78 32
rect -64 -44 -60 41
rect -12 19 68 23
rect -50 -33 -46 -4
rect -12 -13 -8 19
rect 5 -8 11 -3
rect 45 -8 51 -4
rect 5 -33 9 -8
rect -50 -37 9 -33
rect 47 -34 51 -8
rect -64 -78 -61 -49
rect -37 -56 -33 -37
rect 5 -50 9 -37
rect 45 -39 51 -34
rect 5 -55 18 -50
rect -39 -60 -33 -56
rect -29 -78 -25 -62
rect 41 -78 45 -39
rect -64 -82 45 -78
rect 64 -87 68 19
rect -12 -100 77 -96
rect -82 -109 -60 -105
rect -64 -163 -60 -109
rect -50 -152 -46 -123
rect -12 -132 -8 -100
rect 5 -127 11 -122
rect 45 -127 51 -123
rect 5 -152 9 -127
rect -50 -156 9 -152
rect 47 -153 51 -127
rect -64 -197 -61 -168
rect -37 -175 -33 -156
rect 5 -169 9 -156
rect 45 -158 51 -153
rect 5 -174 18 -169
rect -39 -179 -33 -175
rect -29 -197 -25 -181
rect 41 -197 45 -158
rect -64 -201 45 -197
rect 64 -236 68 -109
rect 73 -227 77 -100
rect 89 -105 93 32
rect 107 -44 111 41
rect 159 19 238 23
rect 121 -33 125 -4
rect 159 -13 163 19
rect 176 -8 182 -3
rect 216 -8 222 -4
rect 176 -33 180 -8
rect 121 -37 180 -33
rect 218 -34 222 -8
rect 107 -78 110 -49
rect 134 -56 138 -37
rect 176 -50 180 -37
rect 216 -39 222 -34
rect 176 -55 189 -50
rect 132 -60 138 -56
rect 142 -78 146 -62
rect 212 -78 216 -39
rect 107 -82 216 -78
rect 234 -87 238 19
rect 159 -100 247 -96
rect 89 -109 111 -105
rect 107 -163 111 -109
rect 121 -152 125 -123
rect 159 -132 163 -100
rect 176 -127 182 -122
rect 216 -127 222 -123
rect 176 -152 180 -127
rect 121 -156 180 -152
rect 218 -153 222 -127
rect 107 -197 110 -168
rect 134 -175 138 -156
rect 176 -169 180 -156
rect 216 -158 222 -153
rect 176 -174 189 -169
rect 132 -179 138 -175
rect 142 -197 146 -181
rect 212 -197 216 -158
rect 107 -201 216 -197
rect 234 -236 238 -109
rect 243 -228 247 -100
<< labels >>
rlabel metal1 172 -85 174 -84 1 gnd
rlabel metal1 172 25 174 26 5 vdd
rlabel metal1 172 -94 174 -93 5 vdd
rlabel metal1 172 -204 174 -203 1 gnd
rlabel metal1 1 -85 3 -84 1 gnd
rlabel metal1 1 25 3 26 5 vdd
rlabel metal1 1 -94 3 -93 5 vdd
rlabel metal1 1 -204 3 -203 1 gnd
rlabel ndcontact 27 -186 28 -185 1 xr03
rlabel ndcontact 27 -164 28 -163 1 xr02
rlabel pdcontact 27 -138 28 -137 1 xr01
rlabel pdcontact 27 -116 28 -115 1 xr00
rlabel metal1 -12 -183 -11 -182 1 b0_bar
rlabel metal1 -42 -183 -41 -182 1 a0_bar
rlabel metal1 -68 -166 -66 -165 3 b0
rlabel metal1 -68 -179 -66 -178 3 a0
rlabel pdcontact -32 -113 -31 -111 1 an0
rlabel metal1 -68 -60 -66 -59 1 a1
rlabel metal1 -68 -47 -66 -46 1 b1
rlabel metal1 -43 -64 -41 -63 1 a1_bar
rlabel metal1 -13 -64 -11 -63 1 b1_bar
rlabel pdcontact -32 5 -31 7 1 an1
rlabel pdcontact 27 1 28 3 1 xr10
rlabel pdcontact 27 -21 28 -19 1 xr11
rlabel ndcontact 27 -45 28 -44 1 xr12
rlabel ndcontact 27 -67 28 -66 1 xr13
rlabel metal1 103 -179 105 -178 1 a2
rlabel metal1 103 -166 105 -165 1 b2
rlabel metal1 128 -183 130 -182 1 a2_bar
rlabel pdcontact 139 -114 140 -112 1 an2
rlabel metal1 103 -60 105 -59 1 a3
rlabel metal1 103 -47 105 -46 1 b3
rlabel metal1 128 -64 130 -63 1 a3_bar
rlabel metal1 158 -64 160 -63 1 b3_bar
rlabel pdcontact 139 5 140 7 1 an3
rlabel pdcontact 198 -118 199 -116 1 xr20
rlabel pdcontact 198 -139 199 -137 1 xr21
rlabel ndcontact 198 -164 199 -163 1 xr22
rlabel ndcontact 198 -186 199 -185 1 xr23
rlabel metal1 -90 -213 -88 -212 3 a0
rlabel metal1 -89 -222 -87 -221 3 a1
rlabel metal1 -89 -231 -87 -230 3 a2
rlabel metal1 -89 -240 -87 -239 2 a3
rlabel metal1 -90 -204 -88 -203 3 gnd
rlabel metal1 -89 33 -87 34 3 b0
rlabel metal1 -89 42 -87 43 3 b1
rlabel metal1 -89 51 -87 52 3 b2
rlabel metal1 -89 61 -87 62 4 b3
rlabel metal1 -89 25 -87 26 3 vdd
rlabel pdcontact 198 1 199 3 1 xr30
rlabel pdcontact 198 -21 199 -19 1 xr31
rlabel ndcontact 198 -45 199 -44 1 xr32
rlabel ndcontact 198 -67 199 -66 1 xr33
rlabel metal1 254 -205 256 -204 1 gnd
rlabel metal1 254 -213 256 -212 1 g0
rlabel metal1 254 -222 256 -221 1 g1
rlabel metal1 254 -231 256 -230 1 g2
rlabel metal1 254 -240 256 -239 1 g3
rlabel metal1 258 24 260 25 1 vdd
rlabel metal1 258 33 260 34 1 p0
rlabel metal1 258 42 260 43 1 p1
rlabel metal1 258 50 260 51 1 p2
rlabel metal1 258 60 260 61 5 p3
rlabel metal1 158 -183 160 -182 1 b2_bar
<< end >>
